
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;
use ieee.numeric_std.all;
use work.convolution_pkg.all;

architecture fake_memory_dog of input_ram is
    type memory_assembly is array(0 to padded_dog_size) of std_logic_vector(15 downto 0);
  signal memory : memory_assembly := (
  x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"00AD",
x"00AD",
x"00AA",
x"00AB",
x"00AB",
x"00A9",
x"00AA",
x"00AC",
x"00AA",
x"00A9",
x"00AA",
x"00A8",
x"00A9",
x"00AD",
x"00AE",
x"00AB",
x"00AA",
x"00AD",
x"00AB",
x"00AC",
x"00AC",
x"00AC",
x"00AD",
x"00B0",
x"00AF",
x"00AF",
x"00B0",
x"00B1",
x"00B1",
x"00AF",
x"00B0",
x"00AF",
x"00AF",
x"00B1",
x"00B1",
x"00B1",
x"00B3",
x"00B3",
x"00B1",
x"00B2",
x"00B1",
x"00B2",
x"00B2",
x"00B0",
x"00B0",
x"00B2",
x"00B1",
x"00AD",
x"00AE",
x"00AE",
x"00AE",
x"00AF",
x"00AF",
x"00AE",
x"00AD",
x"00B0",
x"00AE",
x"00AF",
x"00B1",
x"00B0",
x"00B0",
x"00B1",
x"00B1",
x"00B1",
x"00B2",
x"00B3",
x"00B1",
x"00B2",
x"00B1",
x"00B1",
x"00AF",
x"00B2",
x"00AB",
x"0092",
x"0085",
x"0080",
x"007F",
x"0079",
x"008E",
x"008C",
x"0062",
x"0052",
x"0058",
x"007C",
x"007E",
x"007B",
x"007B",
x"0084",
x"007B",
x"0087",
x"009C",
x"009A",
x"009A",
x"009E",
x"009B",
x"0097",
x"0097",
x"0093",
x"0092",
x"0096",
x"0091",
x"0098",
x"0099",
x"009D",
x"0098",
x"008E",
x"0096",
x"008A",
x"0086",
x"008A",
x"008F",
x"0089",
x"008D",
x"008D",
x"008C",
x"0084",
x"0083",
x"008A",
x"009B",
x"0095",
x"008B",
x"0097",
x"0096",
x"0080",
x"0091",
x"0088",
x"008A",
x"008E",
x"0000",
x"0000",
x"0000",
x"0000",
x"00AC",
x"00AC",
x"00AC",
x"00AC",
x"00AC",
x"00AB",
x"00AA",
x"00AE",
x"00AC",
x"00AA",
x"00AB",
x"00AA",
x"00A9",
x"00AA",
x"00AE",
x"00AC",
x"00AC",
x"00AC",
x"00AB",
x"00AA",
x"00AE",
x"00AE",
x"00AE",
x"00B1",
x"00B0",
x"00AF",
x"00B1",
x"00B0",
x"00B0",
x"00B1",
x"00B1",
x"00B0",
x"00AF",
x"00B2",
x"00B2",
x"00B1",
x"00B2",
x"00B3",
x"00B2",
x"00B4",
x"00B1",
x"00B2",
x"00B3",
x"00B3",
x"00B2",
x"00B1",
x"00B0",
x"00AF",
x"00AF",
x"00AE",
x"00AE",
x"00B0",
x"00AE",
x"00AD",
x"00AE",
x"00B0",
x"00B0",
x"00B0",
x"00B1",
x"00B1",
x"00B1",
x"00B0",
x"00B1",
x"00B0",
x"00B1",
x"00B2",
x"00B1",
x"00B2",
x"00B1",
x"00B1",
x"00B2",
x"00B2",
x"00AF",
x"0094",
x"0085",
x"007F",
x"0081",
x"0076",
x"0083",
x"0098",
x"0060",
x"004D",
x"0057",
x"0089",
x"0094",
x"0094",
x"0096",
x"0086",
x"008A",
x"009D",
x"0099",
x"0099",
x"009B",
x"009E",
x"0099",
x"0097",
x"0093",
x"0092",
x"0096",
x"0095",
x"0097",
x"009D",
x"0095",
x"0099",
x"009A",
x"0096",
x"0093",
x"0090",
x"008C",
x"0096",
x"0091",
x"008F",
x"0088",
x"0093",
x"0090",
x"0084",
x"0086",
x"008F",
x"009E",
x"00A4",
x"008E",
x"008D",
x"0081",
x"007F",
x"0087",
x"0080",
x"0080",
x"0093",
x"0000",
x"0000",
x"0000",
x"0000",
x"00AD",
x"00AD",
x"00AC",
x"00AB",
x"00AD",
x"00AB",
x"00AC",
x"00AD",
x"00AB",
x"00AB",
x"00AD",
x"00AB",
x"00AA",
x"00AC",
x"00AC",
x"00AB",
x"00AC",
x"00AE",
x"00AB",
x"00AC",
x"00AF",
x"00AD",
x"00AE",
x"00B1",
x"00B1",
x"00B0",
x"00B0",
x"00B0",
x"00B1",
x"00B2",
x"00B1",
x"00AE",
x"00B0",
x"00B3",
x"00B2",
x"00B1",
x"00B3",
x"00B4",
x"00B4",
x"00B3",
x"00B2",
x"00B2",
x"00B2",
x"00B3",
x"00B1",
x"00B2",
x"00B1",
x"00B0",
x"00B0",
x"00B0",
x"00B0",
x"00B0",
x"00B0",
x"00AE",
x"00AF",
x"00AF",
x"00AF",
x"00AF",
x"00B2",
x"00B1",
x"00B1",
x"00B1",
x"00B2",
x"00B2",
x"00B2",
x"00B1",
x"00AF",
x"00B1",
x"00B1",
x"00B1",
x"00B1",
x"00B2",
x"00AB",
x"0091",
x"0083",
x"0080",
x"0082",
x"0079",
x"0076",
x"007C",
x"005D",
x"004D",
x"0057",
x"0084",
x"0093",
x"00A2",
x"0099",
x"009F",
x"0098",
x"0092",
x"0098",
x"0097",
x"00A3",
x"00A1",
x"009B",
x"0094",
x"0092",
x"0092",
x"0096",
x"009E",
x"0099",
x"009C",
x"009B",
x"009C",
x"0099",
x"0096",
x"0097",
x"008D",
x"0086",
x"0091",
x"008D",
x"008B",
x"0089",
x"009B",
x"0095",
x"008B",
x"007F",
x"008B",
x"0097",
x"00A3",
x"0091",
x"0089",
x"007B",
x"0079",
x"008A",
x"0090",
x"0086",
x"009A",
x"0000",
x"0000",
x"0000",
x"0000",
x"00AD",
x"00AD",
x"00AB",
x"00AB",
x"00AE",
x"00AC",
x"00AD",
x"00AD",
x"00AB",
x"00AA",
x"00AE",
x"00AB",
x"00AB",
x"00AC",
x"00AE",
x"00AE",
x"00AC",
x"00AD",
x"00AE",
x"00AD",
x"00B0",
x"00AE",
x"00AF",
x"00B2",
x"00B1",
x"00AF",
x"00B1",
x"00B2",
x"00B1",
x"00B1",
x"00B0",
x"00AF",
x"00B0",
x"00B3",
x"00B2",
x"00B2",
x"00B3",
x"00B5",
x"00B3",
x"00B4",
x"00B4",
x"00B3",
x"00B3",
x"00B3",
x"00B2",
x"00B1",
x"00B2",
x"00AF",
x"00B1",
x"00B1",
x"00B0",
x"00B0",
x"00B0",
x"00B0",
x"00B1",
x"00B1",
x"00B1",
x"00B0",
x"00B1",
x"00B1",
x"00B1",
x"00B3",
x"00B3",
x"00B2",
x"00B1",
x"00B1",
x"00B0",
x"00B1",
x"00B1",
x"00B1",
x"00B1",
x"00B3",
x"00A6",
x"008C",
x"0087",
x"0083",
x"007F",
x"0070",
x"006B",
x"007B",
x"0060",
x"004D",
x"0055",
x"007A",
x"0089",
x"0095",
x"0092",
x"00BA",
x"00A8",
x"008E",
x"0098",
x"009E",
x"00A3",
x"009E",
x"0098",
x"0094",
x"0092",
x"0092",
x"0095",
x"009A",
x"009C",
x"009D",
x"00A0",
x"009E",
x"0098",
x"0098",
x"009A",
x"008E",
x"007F",
x"0093",
x"008D",
x"0087",
x"0099",
x"009E",
x"008B",
x"0082",
x"0086",
x"008D",
x"0098",
x"00A7",
x"008D",
x"008E",
x"0088",
x"008E",
x"0085",
x"0089",
x"0091",
x"00A4",
x"0000",
x"0000",
x"0000",
x"0000",
x"00AD",
x"00AD",
x"00AC",
x"00AC",
x"00AF",
x"00AC",
x"00AE",
x"00AF",
x"00AD",
x"00AB",
x"00AD",
x"00AD",
x"00AC",
x"00AE",
x"00AE",
x"00AE",
x"00AF",
x"00AF",
x"00AE",
x"00AF",
x"00B1",
x"00B1",
x"00B0",
x"00B2",
x"00B1",
x"00B0",
x"00B3",
x"00B5",
x"00B3",
x"00B3",
x"00B3",
x"00B1",
x"00B1",
x"00B2",
x"00B2",
x"00B3",
x"00B4",
x"00B5",
x"00B4",
x"00B6",
x"00B6",
x"00B6",
x"00B4",
x"00B3",
x"00B2",
x"00B2",
x"00B2",
x"00B0",
x"00B1",
x"00B1",
x"00B1",
x"00B2",
x"00AF",
x"00B0",
x"00B1",
x"00B1",
x"00B1",
x"00B0",
x"00B1",
x"00B1",
x"00B2",
x"00B2",
x"00B2",
x"00B2",
x"00B2",
x"00B1",
x"00B1",
x"00B1",
x"00B1",
x"00B2",
x"00B3",
x"00B2",
x"00A6",
x"008F",
x"0087",
x"0081",
x"007C",
x"007D",
x"00AD",
x"00A6",
x"0068",
x"004A",
x"0055",
x"0080",
x"008E",
x"0093",
x"0096",
x"00B0",
x"00A3",
x"008E",
x"0099",
x"0099",
x"00A1",
x"00A1",
x"0098",
x"0097",
x"0090",
x"0094",
x"0092",
x"0097",
x"009A",
x"009E",
x"009B",
x"0096",
x"0098",
x"009F",
x"009B",
x"0087",
x"0081",
x"0094",
x"008E",
x"008E",
x"009D",
x"009E",
x"008E",
x"007F",
x"007B",
x"0096",
x"00A0",
x"0099",
x"008E",
x"008D",
x"009A",
x"0090",
x"008D",
x"008A",
x"0092",
x"00A6",
x"0000",
x"0000",
x"0000",
x"0000",
x"00AD",
x"00AC",
x"00A9",
x"00AB",
x"00AF",
x"00AE",
x"00AF",
x"00AF",
x"00AC",
x"00AB",
x"00AF",
x"00AD",
x"00AE",
x"00B0",
x"00B0",
x"00AE",
x"00B0",
x"00B1",
x"00AF",
x"00AF",
x"00B1",
x"00B0",
x"00B0",
x"00B3",
x"00B2",
x"00B2",
x"00B4",
x"00B5",
x"00B5",
x"00B4",
x"00B4",
x"00B3",
x"00B3",
x"00B2",
x"00B1",
x"00B3",
x"00B5",
x"00B6",
x"00B5",
x"00B7",
x"00B6",
x"00B5",
x"00B6",
x"00B5",
x"00B1",
x"00B2",
x"00B2",
x"00B0",
x"00B2",
x"00B1",
x"00B2",
x"00B2",
x"00B1",
x"00B1",
x"00B1",
x"00B2",
x"00B1",
x"00B1",
x"00B3",
x"00B3",
x"00B2",
x"00B2",
x"00B1",
x"00B1",
x"00B2",
x"00B2",
x"00B2",
x"00B1",
x"00B2",
x"00B4",
x"00B1",
x"00AE",
x"00A9",
x"0096",
x"0086",
x"007C",
x"0079",
x"0086",
x"00B3",
x"009C",
x"0064",
x"004C",
x"0056",
x"0081",
x"008E",
x"0099",
x"009C",
x"0089",
x"0099",
x"0092",
x"009A",
x"0092",
x"009D",
x"009F",
x"0097",
x"0094",
x"0091",
x"0094",
x"0095",
x"0099",
x"009B",
x"009E",
x"009D",
x"0097",
x"0096",
x"009B",
x"0097",
x"0087",
x"007E",
x"0098",
x"0095",
x"0096",
x"0098",
x"008E",
x"0094",
x"0089",
x"007F",
x"008A",
x"009B",
x"0098",
x"0098",
x"0098",
x"00A5",
x"0090",
x"008E",
x"008F",
x"007B",
x"0092",
x"0000",
x"0000",
x"0000",
x"0000",
x"00AF",
x"00AE",
x"00AC",
x"00AD",
x"00AE",
x"00AE",
x"00AF",
x"00B0",
x"00AD",
x"00AC",
x"00AF",
x"00AE",
x"00AF",
x"00B0",
x"00B0",
x"00B0",
x"00B1",
x"00B2",
x"00AE",
x"00AF",
x"00B0",
x"00B0",
x"00B0",
x"00B3",
x"00B2",
x"00B3",
x"00B5",
x"00B5",
x"00B5",
x"00B6",
x"00B6",
x"00B4",
x"00B4",
x"00B4",
x"00B2",
x"00B3",
x"00B4",
x"00B7",
x"00B5",
x"00B7",
x"00B5",
x"00B4",
x"00B6",
x"00B4",
x"00B2",
x"00B3",
x"00B2",
x"00B2",
x"00B2",
x"00B1",
x"00B2",
x"00B4",
x"00B3",
x"00B1",
x"00B2",
x"00B2",
x"00B1",
x"00B1",
x"00B2",
x"00B3",
x"00B1",
x"00B2",
x"00B1",
x"00B2",
x"00B2",
x"00B1",
x"00B1",
x"00B2",
x"00B2",
x"00B2",
x"00B2",
x"00B2",
x"00B1",
x"0098",
x"0086",
x"0080",
x"0081",
x"0084",
x"00A8",
x"00A8",
x"005C",
x"004E",
x"0059",
x"007F",
x"0087",
x"008E",
x"0091",
x"007D",
x"0097",
x"0096",
x"009A",
x"0097",
x"009F",
x"009E",
x"0097",
x"008F",
x"0092",
x"0095",
x"009A",
x"009C",
x"009E",
x"0099",
x"0098",
x"009A",
x"00A0",
x"00A3",
x"0095",
x"0087",
x"0085",
x"0090",
x"008B",
x"0090",
x"008E",
x"0094",
x"0096",
x"0084",
x"0089",
x"0090",
x"0090",
x"0091",
x"0091",
x"0086",
x"0095",
x"0094",
x"0087",
x"0085",
x"008A",
x"0093",
x"0000",
x"0000",
x"0000",
x"0000",
x"00AF",
x"00AF",
x"00AE",
x"00AE",
x"00AF",
x"00AF",
x"00AF",
x"00B1",
x"00AF",
x"00AF",
x"00B0",
x"00AE",
x"00AE",
x"00B0",
x"00B2",
x"00B2",
x"00B0",
x"00B1",
x"00B0",
x"00B0",
x"00B1",
x"00B1",
x"00B1",
x"00B2",
x"00B5",
x"00B3",
x"00B5",
x"00B6",
x"00B7",
x"00B7",
x"00B5",
x"00B6",
x"00B5",
x"00B5",
x"00B4",
x"00B3",
x"00B5",
x"00B8",
x"00B7",
x"00B6",
x"00B7",
x"00B6",
x"00B6",
x"00B5",
x"00B3",
x"00B3",
x"00B2",
x"00B2",
x"00B2",
x"00B2",
x"00B1",
x"00B3",
x"00B2",
x"00B2",
x"00B2",
x"00B2",
x"00B3",
x"00B2",
x"00B3",
x"00B3",
x"00B0",
x"00B1",
x"00B1",
x"00B0",
x"00B2",
x"00B1",
x"00B1",
x"00B1",
x"00B2",
x"00B2",
x"00B2",
x"00B3",
x"00B3",
x"00A3",
x"0092",
x"0089",
x"008D",
x"008E",
x"00B2",
x"009F",
x"005B",
x"004E",
x"005A",
x"0087",
x"0094",
x"0099",
x"0097",
x"007C",
x"0093",
x"0096",
x"0097",
x"0097",
x"00A3",
x"00A0",
x"0098",
x"0091",
x"008F",
x"0099",
x"009A",
x"00A2",
x"00A2",
x"0099",
x"0097",
x"0095",
x"009B",
x"00A2",
x"009B",
x"0083",
x"0090",
x"009D",
x"0092",
x"0090",
x"0090",
x"009C",
x"008D",
x"0081",
x"0077",
x"0086",
x"008F",
x"008E",
x"0083",
x"0089",
x"008A",
x"0090",
x"008C",
x"0091",
x"0091",
x"0097",
x"0000",
x"0000",
x"0000",
x"0000",
x"00B1",
x"00B0",
x"00AD",
x"00AF",
x"00B0",
x"00AE",
x"00AF",
x"00B1",
x"00B1",
x"00B0",
x"00B1",
x"00B1",
x"00AE",
x"00B2",
x"00B2",
x"00B1",
x"00B1",
x"00B2",
x"00B1",
x"00B2",
x"00B1",
x"00B0",
x"00B2",
x"00B4",
x"00B4",
x"00B3",
x"00B6",
x"00B7",
x"00B6",
x"00B9",
x"00B7",
x"00B5",
x"00B6",
x"00B7",
x"00B6",
x"00B6",
x"00B6",
x"00B6",
x"00B8",
x"00B9",
x"00B7",
x"00B5",
x"00B7",
x"00B7",
x"00B5",
x"00B3",
x"00B2",
x"00B1",
x"00B2",
x"00B2",
x"00B1",
x"00B4",
x"00B2",
x"00B2",
x"00B2",
x"00B3",
x"00B2",
x"00B2",
x"00B3",
x"00B0",
x"00B1",
x"00B2",
x"00B1",
x"00B0",
x"00B2",
x"00B2",
x"00B1",
x"00B1",
x"00B0",
x"00B1",
x"00B1",
x"00B3",
x"00B2",
x"00AA",
x"00A3",
x"0094",
x"0099",
x"008F",
x"00AF",
x"0097",
x"0059",
x"004E",
x"005C",
x"0083",
x"008E",
x"0099",
x"0097",
x"007C",
x"007E",
x"008C",
x"0098",
x"0094",
x"00A2",
x"009F",
x"0097",
x"0090",
x"008D",
x"0098",
x"009C",
x"00A3",
x"00A5",
x"009C",
x"0099",
x"0093",
x"009A",
x"0099",
x"0096",
x"007E",
x"0096",
x"009D",
x"008E",
x"0083",
x"0090",
x"009D",
x"008B",
x"007E",
x"007F",
x"0095",
x"0095",
x"008C",
x"0089",
x"0093",
x"008E",
x"0089",
x"008E",
x"008D",
x"0085",
x"008D",
x"0000",
x"0000",
x"0000",
x"0000",
x"00B0",
x"00AF",
x"00AF",
x"00B0",
x"00B0",
x"00AE",
x"00AF",
x"00B2",
x"00B1",
x"00B2",
x"00B1",
x"00B0",
x"00AE",
x"00B1",
x"00B2",
x"00B1",
x"00B2",
x"00B2",
x"00B2",
x"00B1",
x"00B2",
x"00B0",
x"00B2",
x"00B6",
x"00B4",
x"00B4",
x"00B7",
x"00B6",
x"00B6",
x"00C1",
x"00BB",
x"00B5",
x"00B7",
x"00B8",
x"00B5",
x"00B6",
x"00B7",
x"00B7",
x"00B9",
x"00BA",
x"00B8",
x"00B7",
x"00B6",
x"00B6",
x"00B4",
x"00B4",
x"00B4",
x"00B2",
x"00B3",
x"00B4",
x"00B2",
x"00B5",
x"00B3",
x"00B2",
x"00B1",
x"00B3",
x"00B1",
x"00B3",
x"00B4",
x"00B1",
x"00B1",
x"00B3",
x"00B1",
x"00B1",
x"00B2",
x"00B2",
x"00B1",
x"00B1",
x"00B0",
x"00B2",
x"00B2",
x"00B3",
x"00B1",
x"00B0",
x"00AF",
x"00AD",
x"00AA",
x"0096",
x"00A4",
x"008B",
x"005B",
x"004E",
x"005D",
x"007F",
x"0086",
x"0095",
x"0096",
x"0088",
x"007A",
x"0085",
x"009A",
x"0095",
x"00A0",
x"009F",
x"0093",
x"008E",
x"008E",
x"009B",
x"00A0",
x"00A2",
x"009E",
x"0091",
x"009A",
x"0097",
x"009A",
x"0094",
x"0094",
x"0087",
x"009B",
x"0093",
x"008C",
x"0085",
x"008E",
x"009D",
x"009A",
x"0085",
x"008E",
x"0091",
x"008C",
x"0091",
x"007E",
x"009A",
x"0095",
x"008A",
x"0088",
x"0084",
x"008F",
x"008A",
x"0000",
x"0000",
x"0000",
x"0000",
x"00B1",
x"00B1",
x"00B0",
x"00B0",
x"00AE",
x"00AF",
x"00AF",
x"00B3",
x"00B2",
x"00B0",
x"00B1",
x"00B0",
x"00AF",
x"00B2",
x"00B3",
x"00B3",
x"00B2",
x"00B2",
x"00B1",
x"00B2",
x"00B2",
x"00B2",
x"00B5",
x"00B6",
x"00B5",
x"00B4",
x"00B7",
x"00B7",
x"00B6",
x"00B8",
x"00B9",
x"00B5",
x"00B7",
x"00B8",
x"00B4",
x"00B5",
x"00B7",
x"00B7",
x"00B8",
x"00B9",
x"00B7",
x"00B7",
x"00B7",
x"00B7",
x"00B4",
x"00B5",
x"00B5",
x"00B2",
x"00B2",
x"00B3",
x"00B2",
x"00B4",
x"00B3",
x"00B1",
x"00B2",
x"00B3",
x"00B1",
x"00B2",
x"00B4",
x"00B1",
x"00B0",
x"00B3",
x"00B1",
x"00B2",
x"00B1",
x"00B1",
x"00B2",
x"00B2",
x"00B2",
x"00B2",
x"00B2",
x"00B2",
x"00B1",
x"00B3",
x"00B2",
x"00B2",
x"00AF",
x"00A4",
x"00B5",
x"008F",
x"005D",
x"004E",
x"005D",
x"0087",
x"0091",
x"0096",
x"009F",
x"00AB",
x"009E",
x"0090",
x"0099",
x"0094",
x"00A0",
x"009E",
x"0096",
x"0092",
x"008D",
x"0097",
x"009F",
x"00A0",
x"009B",
x"0094",
x"0094",
x"0094",
x"009D",
x"0099",
x"0098",
x"008F",
x"0096",
x"0097",
x"0094",
x"0093",
x"0090",
x"0097",
x"008C",
x"0086",
x"0098",
x"009B",
x"0095",
x"0092",
x"0088",
x"0096",
x"0089",
x"0094",
x"0099",
x"008A",
x"0083",
x"0091",
x"0000",
x"0000",
x"0000",
x"0000",
x"00B1",
x"00B1",
x"00AF",
x"00AF",
x"00B0",
x"00AF",
x"00B1",
x"00B2",
x"00B0",
x"00B1",
x"00B0",
x"00B0",
x"00B0",
x"00B1",
x"00B2",
x"00B2",
x"00B4",
x"00B4",
x"00B2",
x"00B2",
x"00B2",
x"00B3",
x"00B4",
x"00B7",
x"00B4",
x"00B3",
x"00B7",
x"00B7",
x"00B5",
x"00B7",
x"00B8",
x"00B6",
x"00B7",
x"00B5",
x"00B5",
x"00B6",
x"00B7",
x"00B8",
x"00B8",
x"00B8",
x"00B7",
x"00B6",
x"00B5",
x"00B6",
x"00B5",
x"00B4",
x"00B4",
x"00B2",
x"00B2",
x"00B4",
x"00B2",
x"00B3",
x"00B2",
x"00B1",
x"00B1",
x"00B4",
x"00B2",
x"00B1",
x"00B3",
x"00B2",
x"00B2",
x"00B3",
x"00B2",
x"00B2",
x"00B2",
x"00B2",
x"00B1",
x"00B2",
x"00B2",
x"00B2",
x"00B3",
x"00B2",
x"00B2",
x"00B2",
x"00B2",
x"00B2",
x"00B5",
x"00B8",
x"00A7",
x"0098",
x"005C",
x"004C",
x"005B",
x"0085",
x"008D",
x"0087",
x"0098",
x"00A8",
x"0097",
x"0096",
x"009D",
x"009B",
x"00A9",
x"009F",
x"0089",
x"0083",
x"0092",
x"0092",
x"0099",
x"009F",
x"0098",
x"008F",
x"008E",
x"0097",
x"00A0",
x"00A0",
x"0099",
x"008F",
x"0094",
x"00A1",
x"0093",
x"0094",
x"0093",
x"009B",
x"0085",
x"0080",
x"008C",
x"0097",
x"009D",
x"0088",
x"0088",
x"0095",
x"0089",
x"0081",
x"0096",
x"007D",
x"008E",
x"00A3",
x"0000",
x"0000",
x"0000",
x"0000",
x"00B1",
x"00B1",
x"00AD",
x"00AE",
x"00B0",
x"00AE",
x"00B0",
x"00B2",
x"00B0",
x"00B1",
x"00B1",
x"00B0",
x"00AF",
x"00B1",
x"00B2",
x"00B2",
x"00B5",
x"00B5",
x"00B3",
x"00B4",
x"00B6",
x"00B5",
x"00B4",
x"00B7",
x"00B5",
x"00B5",
x"00B6",
x"00B7",
x"00B7",
x"00B6",
x"00B6",
x"00B6",
x"00B6",
x"00B5",
x"00B5",
x"00B6",
x"00B6",
x"00B7",
x"00B7",
x"00B7",
x"00B7",
x"00B6",
x"00B7",
x"00B7",
x"00B4",
x"00B3",
x"00B3",
x"00B2",
x"00B3",
x"00B3",
x"00B2",
x"00B4",
x"00B2",
x"00B1",
x"00B2",
x"00B3",
x"00B4",
x"00B2",
x"00B3",
x"00B2",
x"00B2",
x"00B2",
x"00B2",
x"00B3",
x"00B3",
x"00B2",
x"00B1",
x"00B1",
x"00B3",
x"00B4",
x"00B3",
x"00B3",
x"00B3",
x"00B4",
x"00B3",
x"00B2",
x"00CD",
x"00C0",
x"007D",
x"0098",
x"0068",
x"004D",
x"005D",
x"0088",
x"0094",
x"0085",
x"0090",
x"00AF",
x"00A1",
x"00A1",
x"00A3",
x"0081",
x"0064",
x"003F",
x"0016",
x"001A",
x"006B",
x"009A",
x"009B",
x"009B",
x"0097",
x"0091",
x"0091",
x"0095",
x"009C",
x"0096",
x"0093",
x"008E",
x"0097",
x"009B",
x"0097",
x"0091",
x"008C",
x"0096",
x"0092",
x"007C",
x"0082",
x"008F",
x"009F",
x"0092",
x"008B",
x"0095",
x"008F",
x"008B",
x"008F",
x"0077",
x"008D",
x"00B0",
x"0000",
x"0000",
x"0000",
x"0000",
x"00B2",
x"00B1",
x"00B0",
x"00B1",
x"00B1",
x"00B0",
x"00B1",
x"00B4",
x"00B0",
x"00AF",
x"00B2",
x"00B0",
x"00AF",
x"00B3",
x"00B3",
x"00B2",
x"00B6",
x"00B6",
x"00B3",
x"00B6",
x"00B7",
x"00B6",
x"00B6",
x"00B8",
x"00B7",
x"00B7",
x"00B8",
x"00B6",
x"00B8",
x"00B9",
x"00B8",
x"00B7",
x"00B7",
x"00B7",
x"00B7",
x"00B7",
x"00B7",
x"00B8",
x"00B8",
x"00B8",
x"00B8",
x"00B7",
x"00B8",
x"00B5",
x"00B5",
x"00B6",
x"00B6",
x"00B4",
x"00B4",
x"00B4",
x"00B3",
x"00B6",
x"00B4",
x"00B3",
x"00B2",
x"00B2",
x"00B3",
x"00B2",
x"00B4",
x"00B2",
x"00B2",
x"00B3",
x"00B1",
x"00B2",
x"00B2",
x"00B2",
x"00B2",
x"00B3",
x"00B4",
x"00B3",
x"00B5",
x"00B5",
x"00B4",
x"00B4",
x"00B3",
x"00B2",
x"00C7",
x"00B0",
x"0063",
x"008D",
x"006B",
x"004D",
x"005C",
x"0086",
x"009E",
x"0092",
x"009F",
x"00A8",
x"0082",
x"0070",
x"0043",
x"0012",
x"0007",
x"0007",
x"0009",
x"0006",
x"0017",
x"0074",
x"009B",
x"009A",
x"0098",
x"0097",
x"0095",
x"009B",
x"0098",
x"0098",
x"0094",
x"0096",
x"009C",
x"009E",
x"0093",
x"008C",
x"0096",
x"00A0",
x"0095",
x"0076",
x"008A",
x"008D",
x"0096",
x"008D",
x"008B",
x"0098",
x"0094",
x"0087",
x"0088",
x"007F",
x"0088",
x"00A4",
x"0000",
x"0000",
x"0000",
x"0000",
x"00B3",
x"00B3",
x"00B1",
x"00B1",
x"00B4",
x"00B1",
x"00B4",
x"00B4",
x"00B1",
x"00B1",
x"00B2",
x"00B0",
x"00B1",
x"00B3",
x"00B3",
x"00B2",
x"00B5",
x"00B6",
x"00B4",
x"00B6",
x"00B8",
x"00B6",
x"00B8",
x"00B8",
x"00B6",
x"00B7",
x"00BA",
x"00B9",
x"00B8",
x"00B9",
x"00BA",
x"00B8",
x"00B7",
x"00B8",
x"00B8",
x"00B8",
x"00B9",
x"00BA",
x"00BB",
x"00B9",
x"00B8",
x"00B7",
x"00B8",
x"00B6",
x"00B6",
x"00B6",
x"00B6",
x"00B5",
x"00B7",
x"00B4",
x"00B4",
x"00B6",
x"00B6",
x"00B6",
x"00B4",
x"00B4",
x"00B3",
x"00B3",
x"00B4",
x"00B3",
x"00B3",
x"00B3",
x"00B1",
x"00B3",
x"00B4",
x"00B3",
x"00B2",
x"00B3",
x"00B2",
x"00B4",
x"00B3",
x"00B3",
x"00B4",
x"00B5",
x"00B5",
x"00B5",
x"00BC",
x"009B",
x"0069",
x"005E",
x"005B",
x"0050",
x"0061",
x"008A",
x"009C",
x"0085",
x"006C",
x"0041",
x"0014",
x"000A",
x"0008",
x"000B",
x"000B",
x"000B",
x"000B",
x"000B",
x"0008",
x"001C",
x"007D",
x"009C",
x"0094",
x"0093",
x"0098",
x"009D",
x"009E",
x"00A3",
x"00A0",
x"0099",
x"009F",
x"009E",
x"0090",
x"008E",
x"0098",
x"009B",
x"0091",
x"0075",
x"0087",
x"0093",
x"0093",
x"0088",
x"0082",
x"0087",
x"0088",
x"007C",
x"008C",
x"0099",
x"009E",
x"009C",
x"0000",
x"0000",
x"0000",
x"0000",
x"00B3",
x"00B3",
x"00B1",
x"00B2",
x"00B4",
x"00B3",
x"00B4",
x"00B5",
x"00B4",
x"00B4",
x"00B4",
x"00B3",
x"00B2",
x"00B3",
x"00B3",
x"00B3",
x"00B7",
x"00B6",
x"00B4",
x"00B6",
x"00B9",
x"00B6",
x"00B7",
x"00BA",
x"00B6",
x"00B8",
x"00B9",
x"00B9",
x"00B8",
x"00B9",
x"00BA",
x"00B9",
x"00BB",
x"00B9",
x"00B8",
x"00BA",
x"00B9",
x"00BA",
x"00BA",
x"00BA",
x"00B7",
x"00B8",
x"00BA",
x"00B8",
x"00B7",
x"00B8",
x"00B6",
x"00B6",
x"00B7",
x"00B6",
x"00B6",
x"00BC",
x"00BD",
x"00B7",
x"00BC",
x"00BA",
x"00B5",
x"00B5",
x"00B5",
x"00B4",
x"00B3",
x"00B3",
x"00B1",
x"00B3",
x"00B3",
x"00B2",
x"00B3",
x"00B3",
x"00B3",
x"00B3",
x"00B2",
x"00B5",
x"00B4",
x"00B4",
x"00B5",
x"00B6",
x"00CC",
x"009D",
x"0070",
x"0056",
x"0058",
x"0056",
x"005E",
x"0065",
x"0044",
x"001D",
x"000D",
x"000B",
x"000D",
x"000E",
x"0010",
x"0011",
x"000E",
x"000C",
x"000C",
x"000C",
x"000B",
x"0006",
x"002E",
x"0091",
x"009E",
x"0098",
x"00A1",
x"009C",
x"009D",
x"00A5",
x"009D",
x"0098",
x"009E",
x"00A3",
x"0099",
x"0098",
x"00A0",
x"00A6",
x"0097",
x"007E",
x"0091",
x"0091",
x"0093",
x"009A",
x"0095",
x"0090",
x"0087",
x"0086",
x"0094",
x"00A6",
x"009A",
x"009F",
x"0000",
x"0000",
x"0000",
x"0000",
x"00B2",
x"00B2",
x"00B1",
x"00B3",
x"00B6",
x"00B5",
x"00B5",
x"00B6",
x"00B6",
x"00B5",
x"00B6",
x"00B4",
x"00B3",
x"00B6",
x"00B5",
x"00B6",
x"00B8",
x"00B7",
x"00B5",
x"00B7",
x"00B8",
x"00B7",
x"00B8",
x"00B9",
x"00B7",
x"00B8",
x"00BA",
x"00BB",
x"00B9",
x"00BA",
x"00BA",
x"00B8",
x"00BA",
x"00B9",
x"00B9",
x"00B9",
x"00BB",
x"00BB",
x"00BA",
x"00BB",
x"00BA",
x"00B9",
x"00BB",
x"00B9",
x"00B7",
x"00B8",
x"00B9",
x"00B9",
x"00B7",
x"00BB",
x"00C0",
x"009D",
x"0062",
x"004B",
x"006B",
x"00A9",
x"00BC",
x"00B6",
x"00B6",
x"00B5",
x"00B5",
x"00B4",
x"00B3",
x"00B3",
x"00B4",
x"00B3",
x"00B2",
x"00B3",
x"00B4",
x"00B3",
x"00B4",
x"00B6",
x"00B5",
x"00B6",
x"00B6",
x"00B7",
x"00D2",
x"00B1",
x"0076",
x"0056",
x"0046",
x"0030",
x"001C",
x"0013",
x"000E",
x"0010",
x"0011",
x"000F",
x"000C",
x"000F",
x"0011",
x"0011",
x"000F",
x"0011",
x"000E",
x"000A",
x"000C",
x"000C",
x"0008",
x"0060",
x"00A3",
x"009F",
x"00A3",
x"009C",
x"00A4",
x"00AE",
x"00A2",
x"009E",
x"00A4",
x"00A8",
x"00A2",
x"00A1",
x"009D",
x"0097",
x"0085",
x"0084",
x"0097",
x"0085",
x"0085",
x"0094",
x"0093",
x"008D",
x"0077",
x"0071",
x"006A",
x"005E",
x"0051",
x"0050",
x"0000",
x"0000",
x"0000",
x"0000",
x"00B2",
x"00B2",
x"00B3",
x"00B5",
x"00B7",
x"00B5",
x"00B6",
x"00B9",
x"00B7",
x"00B6",
x"00B5",
x"00B3",
x"00B2",
x"00B7",
x"00B6",
x"00B6",
x"00B8",
x"00B9",
x"00B7",
x"00B8",
x"00B8",
x"00B7",
x"00B7",
x"00B9",
x"00B9",
x"00B8",
x"00BA",
x"00BB",
x"00B9",
x"00BB",
x"00BA",
x"00B8",
x"00B8",
x"00BA",
x"00BA",
x"00BA",
x"00BB",
x"00BC",
x"00BA",
x"00BB",
x"00BB",
x"00BB",
x"00BB",
x"00B9",
x"00B8",
x"00B9",
x"00BA",
x"00BA",
x"00C0",
x"00B7",
x"0066",
x"001F",
x"0005",
x"0002",
x"0002",
x"0029",
x"008B",
x"00BD",
x"00B7",
x"00B5",
x"00B3",
x"00B5",
x"00B4",
x"00B2",
x"00B3",
x"00B4",
x"00B3",
x"00B3",
x"00B4",
x"00B4",
x"00B5",
x"00B5",
x"00B5",
x"00B7",
x"00B9",
x"00BE",
x"00CA",
x"00AD",
x"0049",
x"001E",
x"000E",
x"000A",
x"000C",
x"000E",
x"000D",
x"000B",
x"000A",
x"000A",
x"0008",
x"000A",
x"000A",
x"000A",
x"000D",
x"000E",
x"000B",
x"000B",
x"000D",
x"000C",
x"0007",
x"0026",
x"0090",
x"0098",
x"0093",
x"007C",
x"007A",
x"0075",
x"0068",
x"0058",
x"0055",
x"0053",
x"004B",
x"0045",
x"003E",
x"0039",
x"0030",
x"0029",
x"002D",
x"0027",
x"0028",
x"002A",
x"002A",
x"0025",
x"0023",
x"0021",
x"001D",
x"001D",
x"001E",
x"001F",
x"0000",
x"0000",
x"0000",
x"0000",
x"00B4",
x"00B4",
x"00B4",
x"00B6",
x"00B8",
x"00B6",
x"00B6",
x"00B8",
x"00B5",
x"00B5",
x"00B6",
x"00B4",
x"00B4",
x"00B7",
x"00B7",
x"00B6",
x"00B7",
x"00B8",
x"00B7",
x"00B8",
x"00B8",
x"00B7",
x"00B8",
x"00BB",
x"00B9",
x"00BA",
x"00BA",
x"00BB",
x"00BB",
x"00BD",
x"00BB",
x"00B9",
x"00BA",
x"00BB",
x"00BA",
x"00BB",
x"00BA",
x"00BB",
x"00BD",
x"00BD",
x"00BA",
x"00BB",
x"00BD",
x"00BB",
x"00BA",
x"00BA",
x"00BA",
x"00C2",
x"00AD",
x"0044",
x"000C",
x"000F",
x"000C",
x"000A",
x"0006",
x"0003",
x"0016",
x"0081",
x"00C0",
x"00B7",
x"00B6",
x"00B6",
x"00B4",
x"00B4",
x"00B4",
x"00B5",
x"00B5",
x"00B5",
x"00B5",
x"00B5",
x"00B7",
x"00B7",
x"00B9",
x"00C3",
x"00BD",
x"008D",
x"004A",
x"001E",
x"0005",
x"0005",
x"0006",
x"0008",
x"0007",
x"0008",
x"000C",
x"000B",
x"0009",
x"000B",
x"000A",
x"000B",
x"000C",
x"000B",
x"000A",
x"000B",
x"000B",
x"000A",
x"000C",
x"000E",
x"000C",
x"000D",
x"0024",
x"0023",
x"001D",
x"0017",
x"001A",
x"0019",
x"0015",
x"0015",
x"0014",
x"0014",
x"0016",
x"0017",
x"0019",
x"001C",
x"0022",
x"0021",
x"0023",
x"0022",
x"0022",
x"0022",
x"0027",
x"0029",
x"0029",
x"002F",
x"0031",
x"0038",
x"0037",
x"0038",
x"0000",
x"0000",
x"0000",
x"0000",
x"00B4",
x"00B4",
x"00B2",
x"00B6",
x"00B7",
x"00B5",
x"00B6",
x"00B8",
x"00B6",
x"00B5",
x"00B7",
x"00B5",
x"00B6",
x"00B8",
x"00B7",
x"00B7",
x"00BA",
x"00B9",
x"00B8",
x"00B9",
x"00B9",
x"00B9",
x"00B9",
x"00BB",
x"00B9",
x"00BB",
x"00BD",
x"00BB",
x"00BA",
x"00BD",
x"00BD",
x"00B9",
x"00BC",
x"00BB",
x"00BA",
x"00BC",
x"00BB",
x"00BC",
x"00BE",
x"00BD",
x"00BA",
x"00BC",
x"00BE",
x"00BD",
x"00BB",
x"00BC",
x"00C4",
x"00A9",
x"0038",
x"000A",
x"0011",
x"0011",
x"000E",
x"000C",
x"0007",
x"0009",
x"0003",
x"0014",
x"0078",
x"00BC",
x"00B9",
x"00B7",
x"00B6",
x"00B5",
x"00B6",
x"00B5",
x"00B5",
x"00B5",
x"00B6",
x"00B8",
x"00BB",
x"00C3",
x"00B7",
x"0083",
x"003D",
x"000E",
x"0001",
x"0004",
x"0007",
x"0007",
x"0009",
x"000A",
x"000A",
x"000C",
x"000C",
x"000C",
x"000B",
x"000B",
x"000A",
x"000B",
x"000B",
x"000C",
x"000A",
x"000A",
x"000C",
x"000A",
x"000C",
x"000C",
x"000C",
x"000B",
x"0008",
x"000D",
x"0011",
x"000C",
x"000A",
x"000E",
x"0012",
x"0018",
x"001A",
x"0019",
x"001B",
x"0020",
x"001F",
x"0020",
x"002D",
x"0033",
x"0036",
x"0034",
x"0030",
x"002A",
x"0021",
x"0020",
x"0021",
x"0026",
x"002B",
x"0032",
x"0039",
x"003D",
x"0000",
x"0000",
x"0000",
x"0000",
x"00B2",
x"00B2",
x"00B5",
x"00B6",
x"00B8",
x"00B4",
x"00B4",
x"00B7",
x"00B6",
x"00B5",
x"00B6",
x"00B5",
x"00B4",
x"00B6",
x"00B7",
x"00B8",
x"00BA",
x"00B9",
x"00BA",
x"00BB",
x"00BB",
x"00BA",
x"00BA",
x"00BC",
x"00BA",
x"00BB",
x"00BC",
x"00BB",
x"00BA",
x"00BC",
x"00BC",
x"00BB",
x"00BC",
x"00BC",
x"00BA",
x"00BB",
x"00BC",
x"00BC",
x"00BC",
x"00BD",
x"00BB",
x"00BC",
x"00BC",
x"00BD",
x"00BC",
x"00C5",
x"00AB",
x"0039",
x"000A",
x"0012",
x"0013",
x"000D",
x"000F",
x"0012",
x"0009",
x"0008",
x"0009",
x"0004",
x"000C",
x"0079",
x"00BE",
x"00B8",
x"00B6",
x"00B6",
x"00B7",
x"00B6",
x"00B6",
x"00B8",
x"00BA",
x"00C2",
x"00C0",
x"0087",
x"0034",
x"0009",
x"0003",
x"0008",
x"000A",
x"000A",
x"000A",
x"000A",
x"000A",
x"000A",
x"000B",
x"000C",
x"000C",
x"000A",
x"000B",
x"000B",
x"000A",
x"000A",
x"000B",
x"000C",
x"000A",
x"000B",
x"000B",
x"000A",
x"000B",
x"000B",
x"000A",
x"000C",
x"000C",
x"0014",
x"0037",
x"003B",
x"002D",
x"001B",
x"0012",
x"0010",
x"0013",
x"0013",
x"0011",
x"0014",
x"0016",
x"0015",
x"0019",
x"0020",
x"0030",
x"003C",
x"0045",
x"0044",
x"003B",
x"002C",
x"001D",
x"0014",
x"0015",
x"0018",
x"001D",
x"0025",
x"0000",
x"0000",
x"0000",
x"0000",
x"00B6",
x"00B6",
x"00B4",
x"00B7",
x"00B7",
x"00B4",
x"00B5",
x"00B8",
x"00B7",
x"00B6",
x"00B6",
x"00B5",
x"00B4",
x"00B6",
x"00B9",
x"00B8",
x"00BB",
x"00BB",
x"00B9",
x"00BA",
x"00BC",
x"00BA",
x"00BA",
x"00BC",
x"00BB",
x"00BC",
x"00BB",
x"00BB",
x"00BC",
x"00BE",
x"00BC",
x"00BA",
x"00BC",
x"00BD",
x"00BA",
x"00BC",
x"00BC",
x"00BC",
x"00BE",
x"00BC",
x"00BB",
x"00BE",
x"00BD",
x"00BE",
x"00C5",
x"00A8",
x"0034",
x"000B",
x"0010",
x"0013",
x"000E",
x"000A",
x"000D",
x"0010",
x"000A",
x"0007",
x"0008",
x"0007",
x"0005",
x"0011",
x"0089",
x"00BF",
x"00B9",
x"00B9",
x"00BC",
x"00BF",
x"00C2",
x"00C2",
x"00BD",
x"008D",
x"003F",
x"000F",
x"0005",
x"000A",
x"0009",
x"000B",
x"000C",
x"000D",
x"000C",
x"000B",
x"000B",
x"000B",
x"000B",
x"000D",
x"000E",
x"000C",
x"000B",
x"000C",
x"000D",
x"000C",
x"000C",
x"000C",
x"000A",
x"000C",
x"000B",
x"000A",
x"000A",
x"000A",
x"000B",
x"000B",
x"000C",
x"000A",
x"0011",
x"0031",
x"0049",
x"004B",
x"0041",
x"002F",
x"0023",
x"001F",
x"001E",
x"001C",
x"0019",
x"0016",
x"0012",
x"000F",
x"0014",
x"001D",
x"002E",
x"0041",
x"004C",
x"004B",
x"0041",
x"0037",
x"002A",
x"001F",
x"0016",
x"0014",
x"0000",
x"0000",
x"0000",
x"0000",
x"00B7",
x"00B7",
x"00B5",
x"00B7",
x"00B7",
x"00B4",
x"00B6",
x"00B8",
x"00B6",
x"00B6",
x"00B7",
x"00B4",
x"00B4",
x"00B8",
x"00B8",
x"00B8",
x"00BB",
x"00BC",
x"00BA",
x"00BA",
x"00BC",
x"00BB",
x"00BA",
x"00BC",
x"00BB",
x"00BD",
x"00BD",
x"00BA",
x"00BB",
x"00BE",
x"00BD",
x"00BB",
x"00BC",
x"00BC",
x"00BB",
x"00BD",
x"00BC",
x"00BC",
x"00BF",
x"00BE",
x"00BD",
x"00BD",
x"00BF",
x"00C5",
x"00AD",
x"0033",
x"000C",
x"0013",
x"0014",
x"0010",
x"000A",
x"0008",
x"000E",
x"0010",
x"000A",
x"0007",
x"0006",
x"0007",
x"0008",
x"0004",
x"001C",
x"00A1",
x"00C3",
x"00BB",
x"00AD",
x"0089",
x"0067",
x"0052",
x"0033",
x"0012",
x"0009",
x"000D",
x"000C",
x"000C",
x"0008",
x"000A",
x"000C",
x"000D",
x"000B",
x"000C",
x"000C",
x"000E",
x"000E",
x"000F",
x"000E",
x"000D",
x"000B",
x"000B",
x"000D",
x"000D",
x"000F",
x"000E",
x"000B",
x"000B",
x"000C",
x"000B",
x"000B",
x"000B",
x"000A",
x"000B",
x"000C",
x"000E",
x"0007",
x"0006",
x"0013",
x"0032",
x"0049",
x"0049",
x"0044",
x"003E",
x"003A",
x"003A",
x"0035",
x"002E",
x"0028",
x"001F",
x"001C",
x"0015",
x"0011",
x"0018",
x"0029",
x"003E",
x"0047",
x"004A",
x"004C",
x"0042",
x"002F",
x"0026",
x"0000",
x"0000",
x"0000",
x"0000",
x"00B7",
x"00B7",
x"00B5",
x"00B8",
x"00B9",
x"00B7",
x"00B8",
x"00B7",
x"00B7",
x"00B7",
x"00B9",
x"00B7",
x"00B7",
x"00BA",
x"00B9",
x"00B8",
x"00B9",
x"00BC",
x"00BB",
x"00BD",
x"00BD",
x"00BC",
x"00BA",
x"00BB",
x"00BC",
x"00BE",
x"00BC",
x"00BB",
x"00BB",
x"00BF",
x"00BD",
x"00BA",
x"00BD",
x"00BD",
x"00BC",
x"00BD",
x"00BD",
x"00BF",
x"00C1",
x"00C0",
x"00BF",
x"00C0",
x"00C7",
x"00B8",
x"003C",
x"000B",
x"0012",
x"0012",
x"0016",
x"000E",
x"000B",
x"0009",
x"0011",
x"0010",
x"000F",
x"000D",
x"0007",
x"0007",
x"0008",
x"0009",
x"0002",
x"002D",
x"0047",
x"0029",
x"001A",
x"000B",
x"0001",
x"0000",
x"0003",
x"0008",
x"000E",
x"000E",
x"000B",
x"000C",
x"0008",
x"0009",
x"000B",
x"000C",
x"000B",
x"000B",
x"000F",
x"0010",
x"000F",
x"0010",
x"000F",
x"000F",
x"000E",
x"000B",
x"000C",
x"000E",
x"000F",
x"000E",
x"000D",
x"000E",
x"000C",
x"000C",
x"000C",
x"000C",
x"000A",
x"000A",
x"000B",
x"000F",
x"000B",
x"0007",
x"0006",
x"000B",
x"0026",
x"0043",
x"004A",
x"004A",
x"004A",
x"0049",
x"0049",
x"0048",
x"0048",
x"0040",
x"0041",
x"0039",
x"002E",
x"001F",
x"0015",
x"001B",
x"002B",
x"0034",
x"003D",
x"0047",
x"003E",
x"0033",
x"0000",
x"0000",
x"0000",
x"0000",
x"00B7",
x"00B7",
x"00B5",
x"00B8",
x"00B9",
x"00B8",
x"00B9",
x"00B9",
x"00B9",
x"00B8",
x"00BA",
x"00B8",
x"00B7",
x"00BA",
x"00B9",
x"00B9",
x"00BA",
x"00BC",
x"00BB",
x"00BE",
x"00BD",
x"00BC",
x"00BD",
x"00BD",
x"00BC",
x"00BE",
x"00BD",
x"00BE",
x"00BE",
x"00BE",
x"00BB",
x"00BB",
x"00BE",
x"00BE",
x"00BD",
x"00BE",
x"00BE",
x"00BF",
x"00C0",
x"00C1",
x"00C0",
x"00C5",
x"00C3",
x"0054",
x"000A",
x"0011",
x"0013",
x"0013",
x"0015",
x"000B",
x"000E",
x"000B",
x"0013",
x"000E",
x"000D",
x"0012",
x"000A",
x"0008",
x"0009",
x"000A",
x"0008",
x"0003",
x"0003",
x"0003",
x"0005",
x"0006",
x"0006",
x"0006",
x"0008",
x"000B",
x"000C",
x"0011",
x"000D",
x"000C",
x"000B",
x"0009",
x"000B",
x"000B",
x"000C",
x"000B",
x"000D",
x"0010",
x"0010",
x"000F",
x"0012",
x"0011",
x"0010",
x"000C",
x"000E",
x"0010",
x"0010",
x"0010",
x"000E",
x"0010",
x"000E",
x"000C",
x"000D",
x"000E",
x"000C",
x"000B",
x"000D",
x"000F",
x"000D",
x"0009",
x"0009",
x"000C",
x"000A",
x"0022",
x"003B",
x"0043",
x"004A",
x"004B",
x"004B",
x"004E",
x"004E",
x"0049",
x"0051",
x"004E",
x"004A",
x"0046",
x"0038",
x"002B",
x"002D",
x"0032",
x"0033",
x"0038",
x"003A",
x"003D",
x"0000",
x"0000",
x"0000",
x"0000",
x"00B8",
x"00B7",
x"00B6",
x"00B9",
x"00B9",
x"00B6",
x"00B8",
x"00BA",
x"00BA",
x"00BA",
x"00BA",
x"00B8",
x"00B7",
x"00BB",
x"00BA",
x"00B9",
x"00BC",
x"00BE",
x"00BB",
x"00BD",
x"00BD",
x"00BB",
x"00BD",
x"00BE",
x"00BD",
x"00BD",
x"00BD",
x"00BD",
x"00BE",
x"00BE",
x"00BE",
x"00BE",
x"00BF",
x"00BD",
x"00BC",
x"00BE",
x"00BE",
x"00C0",
x"00C0",
x"00C0",
x"00C1",
x"00C7",
x"0065",
x"000E",
x"000E",
x"000F",
x"0014",
x"0015",
x"0015",
x"000B",
x"000B",
x"000D",
x"0012",
x"000C",
x"000D",
x"0014",
x"000D",
x"0008",
x"0009",
x"000A",
x"0009",
x"0008",
x"0008",
x"0007",
x"0009",
x"0008",
x"0008",
x"0006",
x"0008",
x"000B",
x"000B",
x"0010",
x"0010",
x"000E",
x"000E",
x"0009",
x"000B",
x"000B",
x"000A",
x"000A",
x"000C",
x"000E",
x"000F",
x"0010",
x"0010",
x"0010",
x"0010",
x"000C",
x"000D",
x"000E",
x"0010",
x"0010",
x"000F",
x"0010",
x"000D",
x"000D",
x"000D",
x"000F",
x"000D",
x"000C",
x"000E",
x"000F",
x"0011",
x"000A",
x"0009",
x"0009",
x"0007",
x"000C",
x"0022",
x"003A",
x"0048",
x"004B",
x"0046",
x"003E",
x"0040",
x"003E",
x"0040",
x"003E",
x"0039",
x"0037",
x"0032",
x"002F",
x"003C",
x"003C",
x"004B",
x"0056",
x"0048",
x"0042",
x"0000",
x"0000",
x"0000",
x"0000",
x"00B7",
x"00B7",
x"00B7",
x"00B9",
x"00B9",
x"00B7",
x"00B9",
x"00BB",
x"00BA",
x"00BA",
x"00BB",
x"00B9",
x"00B7",
x"00BA",
x"00BB",
x"00BB",
x"00BC",
x"00BE",
x"00BC",
x"00BD",
x"00BF",
x"00BD",
x"00BE",
x"00BF",
x"00BE",
x"00BE",
x"00BF",
x"00BC",
x"00BD",
x"00BF",
x"00BF",
x"00C0",
x"00C0",
x"00BF",
x"00BD",
x"00BF",
x"00BF",
x"00C0",
x"00C2",
x"00C3",
x"00CC",
x"007D",
x"0012",
x"0010",
x"0012",
x"000F",
x"0013",
x"0015",
x"0015",
x"000C",
x"000A",
x"0012",
x"0011",
x"000B",
x"000E",
x"0014",
x"000D",
x"0008",
x"000A",
x"000B",
x"000A",
x"0008",
x"0009",
x"0009",
x"0009",
x"0008",
x"0008",
x"0006",
x"0009",
x"000C",
x"000B",
x"000D",
x"0013",
x"0010",
x"000F",
x"0009",
x"000D",
x"000D",
x"000A",
x"000A",
x"000B",
x"000D",
x"000F",
x"0010",
x"0010",
x"0010",
x"000F",
x"000B",
x"000B",
x"000E",
x"000F",
x"0011",
x"000E",
x"000E",
x"000C",
x"000C",
x"000E",
x"000E",
x"000D",
x"000F",
x"000F",
x"0010",
x"0012",
x"000C",
x"0008",
x"000A",
x"0009",
x"0008",
x"0014",
x"002C",
x"003F",
x"0044",
x"0047",
x"003B",
x"0033",
x"0031",
x"0033",
x"0033",
x"0030",
x"002D",
x"002A",
x"0030",
x"0058",
x"0075",
x"0095",
x"009B",
x"0084",
x"0074",
x"0000",
x"0000",
x"0000",
x"0000",
x"00B8",
x"00B8",
x"00B7",
x"00B9",
x"00B8",
x"00B8",
x"00B9",
x"00BA",
x"00B9",
x"00BB",
x"00BC",
x"00B8",
x"00B9",
x"00BC",
x"00BC",
x"00BC",
x"00BF",
x"00BE",
x"00BD",
x"00BE",
x"00BE",
x"00BD",
x"00BD",
x"00BF",
x"00BF",
x"00C0",
x"00BF",
x"00BF",
x"00C1",
x"00C0",
x"00BE",
x"00BF",
x"00C0",
x"00BE",
x"00BF",
x"00C1",
x"00C0",
x"00C1",
x"00C1",
x"00CB",
x"00A9",
x"0029",
x"000B",
x"000F",
x"0013",
x"0012",
x"0014",
x"0015",
x"0013",
x"000E",
x"000C",
x"0010",
x"000C",
x"000C",
x"0010",
x"0014",
x"000D",
x"0008",
x"000A",
x"000B",
x"0009",
x"0007",
x"0008",
x"000A",
x"0009",
x"0008",
x"0008",
x"0008",
x"0008",
x"000D",
x"000C",
x"000D",
x"0011",
x"0013",
x"0012",
x"000A",
x"000C",
x"0010",
x"000D",
x"000B",
x"000C",
x"000E",
x"000F",
x"0010",
x"0011",
x"000F",
x"000D",
x"000D",
x"000B",
x"000C",
x"000E",
x"000F",
x"000D",
x"000F",
x"000B",
x"000C",
x"000C",
x"000B",
x"000C",
x"000E",
x"0010",
x"0011",
x"0012",
x"000D",
x"0006",
x"0008",
x"0009",
x"0009",
x"000A",
x"001C",
x"0033",
x"0049",
x"004A",
x"0046",
x"0033",
x"002D",
x"0032",
x"0036",
x"0049",
x"0060",
x"0079",
x"008B",
x"0093",
x"0096",
x"0092",
x"0086",
x"0077",
x"0089",
x"0000",
x"0000",
x"0000",
x"0000",
x"00B8",
x"00B8",
x"00B6",
x"00BA",
x"00BB",
x"00B7",
x"00B9",
x"00BA",
x"00B9",
x"00BB",
x"00BD",
x"00B9",
x"00B8",
x"00BB",
x"00B9",
x"00BB",
x"00BE",
x"00BD",
x"00BC",
x"00BF",
x"00BE",
x"00BC",
x"00BE",
x"00C0",
x"00BE",
x"00C0",
x"00BF",
x"00BE",
x"00C0",
x"00C1",
x"00BE",
x"00BE",
x"00BF",
x"00BE",
x"00BE",
x"00C0",
x"00C0",
x"00C3",
x"00C9",
x"00BD",
x"0044",
x"000C",
x"000E",
x"000A",
x"000F",
x"0012",
x"0013",
x"0014",
x"0013",
x"000E",
x"000C",
x"000F",
x"000D",
x"000C",
x"0012",
x"0013",
x"000C",
x"0009",
x"000A",
x"000A",
x"0008",
x"0007",
x"0007",
x"0009",
x"0009",
x"0007",
x"0007",
x"0007",
x"0007",
x"000B",
x"000B",
x"000C",
x"000F",
x"0012",
x"0012",
x"000D",
x"0008",
x"000F",
x"000E",
x"000B",
x"000D",
x"000E",
x"000E",
x"0010",
x"0010",
x"000C",
x"000F",
x"0010",
x"000B",
x"000B",
x"000E",
x"000E",
x"000B",
x"0010",
x"000D",
x"000D",
x"000D",
x"000C",
x"000D",
x"0010",
x"0011",
x"0011",
x"0012",
x"0010",
x"0007",
x"0008",
x"0008",
x"0008",
x"0009",
x"000D",
x"0029",
x"004A",
x"004C",
x"004D",
x"005E",
x"0074",
x"0090",
x"009C",
x"008F",
x"008F",
x"009A",
x"009B",
x"0097",
x"009E",
x"00A4",
x"007F",
x"007A",
x"0089",
x"0000",
x"0000",
x"0000",
x"0000",
x"00B8",
x"00B8",
x"00B7",
x"00BA",
x"00BA",
x"00B9",
x"00BA",
x"00BA",
x"00B9",
x"00BC",
x"00BC",
x"00B9",
x"00B8",
x"00BA",
x"00BA",
x"00BB",
x"00BF",
x"00BD",
x"00BC",
x"00BE",
x"00BE",
x"00BC",
x"00BE",
x"00C0",
x"00BF",
x"00BF",
x"00C1",
x"00BF",
x"00BF",
x"00C1",
x"00C0",
x"00BF",
x"00BF",
x"00BF",
x"00C0",
x"00C0",
x"00C1",
x"00CA",
x"00BC",
x"004D",
x"000C",
x"0012",
x"000D",
x"0009",
x"000A",
x"0010",
x"0015",
x"0015",
x"0013",
x"000F",
x"000A",
x"0008",
x"000B",
x"000D",
x"0012",
x"0013",
x"000C",
x"000A",
x"000A",
x"0009",
x"0007",
x"0007",
x"0007",
x"0009",
x"000B",
x"0007",
x"0006",
x"0006",
x"0006",
x"0009",
x"000D",
x"000C",
x"000F",
x"0010",
x"0013",
x"0011",
x"0007",
x"000B",
x"000E",
x"000B",
x"000D",
x"0010",
x"0010",
x"0010",
x"0010",
x"000D",
x"000F",
x"0012",
x"000D",
x"000B",
x"000B",
x"000D",
x"000C",
x"000F",
x"000E",
x"000F",
x"0010",
x"000F",
x"000F",
x"0011",
x"0012",
x"0012",
x"0010",
x"0013",
x"000B",
x"0007",
x"0007",
x"0006",
x"0008",
x"0009",
x"0018",
x"0043",
x"005E",
x"0088",
x"0090",
x"008B",
x"009D",
x"009E",
x"00AD",
x"009B",
x"009B",
x"009B",
x"00A2",
x"009A",
x"0092",
x"0088",
x"0092",
x"009C",
x"0000",
x"0000",
x"0000",
x"0000",
x"00B8",
x"00B8",
x"00B6",
x"00B9",
x"00BA",
x"00B8",
x"00BB",
x"00BA",
x"00BA",
x"00BD",
x"00BD",
x"00B9",
x"00B8",
x"00BA",
x"00BA",
x"00BA",
x"00BD",
x"00BC",
x"00BC",
x"00C0",
x"00BD",
x"00BD",
x"00BE",
x"00BE",
x"00BE",
x"00C0",
x"00C5",
x"00C1",
x"00BF",
x"00C2",
x"00BF",
x"00BF",
x"00C0",
x"00C0",
x"00C0",
x"00C1",
x"00C9",
x"00BE",
x"004D",
x"000A",
x"0010",
x"0013",
x"000F",
x"000B",
x"0009",
x"000F",
x"0015",
x"0015",
x"000F",
x"000D",
x"000B",
x"0008",
x"0008",
x"0010",
x"0013",
x"0011",
x"000D",
x"000C",
x"000B",
x"0009",
x"0008",
x"0008",
x"0007",
x"0009",
x"000B",
x"0007",
x"0005",
x"0005",
x"0006",
x"0007",
x"000C",
x"000C",
x"000D",
x"0010",
x"0011",
x"0012",
x"000A",
x"0009",
x"000C",
x"000B",
x"000D",
x"0010",
x"0010",
x"000F",
x"000F",
x"000E",
x"000D",
x"0010",
x"000E",
x"000B",
x"000B",
x"000E",
x"000D",
x"000F",
x"0011",
x"0010",
x"0011",
x"0010",
x"000F",
x"0011",
x"0014",
x"0013",
x"0010",
x"0015",
x"0010",
x"0007",
x"0006",
x"0006",
x"0007",
x"0008",
x"0009",
x"001E",
x"002C",
x"0023",
x"002F",
x"0031",
x"0034",
x"003F",
x"004C",
x"004F",
x"005B",
x"0065",
x"006A",
x"006B",
x"006E",
x"006A",
x"0077",
x"007B",
x"0000",
x"0000",
x"0000",
x"0000",
x"00BA",
x"00B8",
x"00B8",
x"00BB",
x"00BD",
x"00BA",
x"00BC",
x"00BD",
x"00BC",
x"00BC",
x"00BC",
x"00B9",
x"00B9",
x"00BA",
x"00BB",
x"00BA",
x"00BD",
x"00BD",
x"00BE",
x"00BF",
x"00BE",
x"00BE",
x"00BE",
x"00BF",
x"00BD",
x"00C0",
x"00C0",
x"00C0",
x"00C0",
x"00C1",
x"00BF",
x"00BE",
x"00C1",
x"00C1",
x"00C2",
x"00CC",
x"00B6",
x"004E",
x"000D",
x"0011",
x"0010",
x"0012",
x"0011",
x"0010",
x"000B",
x"000A",
x"0012",
x"0014",
x"000D",
x"000C",
x"000C",
x"0009",
x"0007",
x"0008",
x"000D",
x"000F",
x"000F",
x"0010",
x"000E",
x"0009",
x"0009",
x"0009",
x"0007",
x"0008",
x"000C",
x"0008",
x"0006",
x"0006",
x"0006",
x"0006",
x"0009",
x"000C",
x"000D",
x"000D",
x"000F",
x"0010",
x"000E",
x"0008",
x"000C",
x"000C",
x"000D",
x"000F",
x"000E",
x"000D",
x"000F",
x"000D",
x"0011",
x"0011",
x"0010",
x"0011",
x"000D",
x"000F",
x"0010",
x"0011",
x"0010",
x"0010",
x"0012",
x"0012",
x"0011",
x"0012",
x"0014",
x"0014",
x"0013",
x"0014",
x"0013",
x"0008",
x"0006",
x"0006",
x"0007",
x"0008",
x"0007",
x"0006",
x"0003",
x"0009",
x"001E",
x"001F",
x"0025",
x"0028",
x"002A",
x"002F",
x"0030",
x"003B",
x"002F",
x"001A",
x"000F",
x"000E",
x"000F",
x"0011",
x"0000",
x"0000",
x"0000",
x"0000",
x"00BA",
x"00BA",
x"00BA",
x"00BE",
x"00BC",
x"00B9",
x"00BC",
x"00BE",
x"00BE",
x"00BE",
x"00BD",
x"00BB",
x"00BA",
x"00BA",
x"00B9",
x"00BB",
x"00BD",
x"00BE",
x"00BF",
x"00C0",
x"00BF",
x"00BE",
x"00BE",
x"00C0",
x"00BD",
x"00C0",
x"00C1",
x"00C0",
x"00C1",
x"00C2",
x"00C0",
x"00BF",
x"00C2",
x"00C7",
x"00C6",
x"0088",
x"0033",
x"0010",
x"0012",
x"0014",
x"0014",
x"0013",
x"000E",
x"000F",
x"0012",
x"000C",
x"000E",
x"0012",
x"000E",
x"000A",
x"000E",
x"000B",
x"0006",
x"0008",
x"000F",
x"0010",
x"000F",
x"0012",
x"0011",
x"0008",
x"0008",
x"000A",
x"0007",
x"0008",
x"000F",
x"000B",
x"0007",
x"0006",
x"0007",
x"0008",
x"0008",
x"000D",
x"000D",
x"000F",
x"0010",
x"0010",
x"0011",
x"000A",
x"0009",
x"000B",
x"000A",
x"000D",
x"000E",
x"000E",
x"000E",
x"000E",
x"000F",
x"0010",
x"000E",
x"000F",
x"000F",
x"0010",
x"0010",
x"0011",
x"0010",
x"0011",
x"0011",
x"0012",
x"0011",
x"0013",
x"0014",
x"0014",
x"0013",
x"0014",
x"0013",
x"000C",
x"0007",
x"0008",
x"0008",
x"0008",
x"0007",
x"0009",
x"0007",
x"000D",
x"0019",
x"001A",
x"002A",
x"003D",
x"0040",
x"0043",
x"0038",
x"004C",
x"0058",
x"0052",
x"0039",
x"0018",
x"000C",
x"0009",
x"0000",
x"0000",
x"0000",
x"0000",
x"00BB",
x"00BC",
x"00BB",
x"00BE",
x"00BC",
x"00B9",
x"00BC",
x"00BC",
x"00BC",
x"00BE",
x"00BD",
x"00BA",
x"00BA",
x"00BB",
x"00BA",
x"00BD",
x"00BE",
x"00BF",
x"00BF",
x"00C1",
x"00C0",
x"00BD",
x"00C0",
x"00C0",
x"00BF",
x"00C1",
x"00C2",
x"00BF",
x"00C1",
x"00C2",
x"00C0",
x"00C0",
x"00C5",
x"00C1",
x"005A",
x"000E",
x"000D",
x"0014",
x"0013",
x"0012",
x"0013",
x"0014",
x"000E",
x"000B",
x"000F",
x"0010",
x"0011",
x"0011",
x"000E",
x"000C",
x"0010",
x"000A",
x"0008",
x"000A",
x"000E",
x"0011",
x"0012",
x"0014",
x"0017",
x"000F",
x"0007",
x"000A",
x"0008",
x"0009",
x"0010",
x"000D",
x"0008",
x"0006",
x"0008",
x"0008",
x"0008",
x"000C",
x"000D",
x"000E",
x"000F",
x"000D",
x"000F",
x"000C",
x"0008",
x"000B",
x"000C",
x"000C",
x"000D",
x"000E",
x"000C",
x"000E",
x"000F",
x"0010",
x"000F",
x"0010",
x"0011",
x"0010",
x"0011",
x"0012",
x"0011",
x"0013",
x"0013",
x"0012",
x"0010",
x"0012",
x"0011",
x"0011",
x"0011",
x"0012",
x"0014",
x"0010",
x"0008",
x"0008",
x"0008",
x"0008",
x"0007",
x"0009",
x"0009",
x"0008",
x"0007",
x"0005",
x"001A",
x"0032",
x"002E",
x"0030",
x"002D",
x"0045",
x"0051",
x"0058",
x"0055",
x"0041",
x"0028",
x"001D",
x"0000",
x"0000",
x"0000",
x"0000",
x"00BD",
x"00BD",
x"00BC",
x"00BE",
x"00BC",
x"00BA",
x"00BB",
x"00BB",
x"00BB",
x"00BF",
x"00BF",
x"00BA",
x"00BB",
x"00BC",
x"00BA",
x"00BE",
x"00C0",
x"00BF",
x"00BE",
x"00C1",
x"00C1",
x"00BF",
x"00BF",
x"00C0",
x"00C0",
x"00C3",
x"00C3",
x"00C0",
x"00C2",
x"00C2",
x"00C1",
x"00C2",
x"00CB",
x"0082",
x"0007",
x"000D",
x"000C",
x"0011",
x"0014",
x"0012",
x"0010",
x"0013",
x"0010",
x"000B",
x"000A",
x"000B",
x"000E",
x"000E",
x"000C",
x"000A",
x"000D",
x"000B",
x"000B",
x"000B",
x"000C",
x"0013",
x"0014",
x"0011",
x"001F",
x"0016",
x"000A",
x"0009",
x"0009",
x"0009",
x"000F",
x"000D",
x"0009",
x"0006",
x"0008",
x"0007",
x"0008",
x"000A",
x"000B",
x"000C",
x"0010",
x"000E",
x"000D",
x"0010",
x"0009",
x"000B",
x"000D",
x"000D",
x"000B",
x"000E",
x"000E",
x"000D",
x"0010",
x"0012",
x"0011",
x"0012",
x"0013",
x"0012",
x"0012",
x"0013",
x"0010",
x"0011",
x"0013",
x"0011",
x"0010",
x"0010",
x"0010",
x"0010",
x"000E",
x"000E",
x"0010",
x"0012",
x"0008",
x"0007",
x"0009",
x"0008",
x"0009",
x"000A",
x"0008",
x"0008",
x"0010",
x"0026",
x"0021",
x"0020",
x"0025",
x"001D",
x"001A",
x"003D",
x"0053",
x"004F",
x"0050",
x"004D",
x"0045",
x"0039",
x"0000",
x"0000",
x"0000",
x"0000",
x"00BF",
x"00BF",
x"00BE",
x"00BE",
x"00BD",
x"00BB",
x"00BB",
x"00BC",
x"00BE",
x"00BF",
x"00BF",
x"00BC",
x"00BC",
x"00BE",
x"00BB",
x"00BD",
x"00BF",
x"00BF",
x"00BD",
x"00C1",
x"00C3",
x"00BF",
x"00C0",
x"00C1",
x"00C2",
x"00C4",
x"00C4",
x"00C0",
x"00C1",
x"00C2",
x"00C2",
x"00C3",
x"00C8",
x"0059",
x"0008",
x"000F",
x"000E",
x"000E",
x"0010",
x"0010",
x"000E",
x"0012",
x"000E",
x"000C",
x"000B",
x"000A",
x"000B",
x"000A",
x"0008",
x"0007",
x"000C",
x"000D",
x"000B",
x"000D",
x"000B",
x"0011",
x"0016",
x"0011",
x"0010",
x"0010",
x"0011",
x"0008",
x"0008",
x"000C",
x"000F",
x"000F",
x"000B",
x"0006",
x"0007",
x"0007",
x"000B",
x"000C",
x"000C",
x"000B",
x"0011",
x"0011",
x"000D",
x"000D",
x"000C",
x"000D",
x"000F",
x"0010",
x"000E",
x"000F",
x"0011",
x"0012",
x"0013",
x"0013",
x"0012",
x"0013",
x"0012",
x"0012",
x"0011",
x"0012",
x"0010",
x"000F",
x"000F",
x"000E",
x"000E",
x"000D",
x"000D",
x"000D",
x"000E",
x"000F",
x"0012",
x"0012",
x"000C",
x"0007",
x"0009",
x"000A",
x"000A",
x"000A",
x"0009",
x"0007",
x"0019",
x"0039",
x"0039",
x"0021",
x"001F",
x"001C",
x"0017",
x"002F",
x"0051",
x"004C",
x"004E",
x"0047",
x"0058",
x"0056",
x"0000",
x"0000",
x"0000",
x"0000",
x"00BF",
x"00BF",
x"00BE",
x"00C0",
x"00BF",
x"00BB",
x"00BD",
x"00BD",
x"00BD",
x"00BF",
x"00BE",
x"00BB",
x"00BB",
x"00BD",
x"00BB",
x"00BC",
x"00BF",
x"00BE",
x"00BF",
x"00C0",
x"00C1",
x"00BF",
x"00C0",
x"00C1",
x"00BF",
x"00C1",
x"00C4",
x"00C1",
x"00C1",
x"00C4",
x"00C2",
x"00C4",
x"00C5",
x"0045",
x"000F",
x"0010",
x"0010",
x"0011",
x"000E",
x"000F",
x"000E",
x"0010",
x"000E",
x"000B",
x"000B",
x"000A",
x"000B",
x"000A",
x"000A",
x"000B",
x"000C",
x"000F",
x"000C",
x"000C",
x"000A",
x"000C",
x"0015",
x"0014",
x"0013",
x"000F",
x"0011",
x"000A",
x"0009",
x"000D",
x"000F",
x"000F",
x"000C",
x"0009",
x"0006",
x"000A",
x"0010",
x"0010",
x"000D",
x"000C",
x"000E",
x"000E",
x"000D",
x"0010",
x"000F",
x"0010",
x"0011",
x"0013",
x"0011",
x"0011",
x"000F",
x"0011",
x"0013",
x"0012",
x"000E",
x"000F",
x"0010",
x"0010",
x"0010",
x"0010",
x"0010",
x"0010",
x"000F",
x"000D",
x"000C",
x"000C",
x"000C",
x"000C",
x"000B",
x"000B",
x"000A",
x"000C",
x"000B",
x"0007",
x"0008",
x"0009",
x"0009",
x"000A",
x"0009",
x"0014",
x"0014",
x"001A",
x"002D",
x"0034",
x"0026",
x"001B",
x"0015",
x"0023",
x"004C",
x"0051",
x"003E",
x"003E",
x"0055",
x"0054",
x"0000",
x"0000",
x"0000",
x"0000",
x"00C1",
x"00C0",
x"00BF",
x"00BF",
x"00BE",
x"00BC",
x"00BE",
x"00BE",
x"00BE",
x"00C0",
x"00C0",
x"00BD",
x"00BB",
x"00BC",
x"00BC",
x"00BD",
x"00BF",
x"00BF",
x"00BE",
x"00C1",
x"00BF",
x"00BE",
x"00BF",
x"00C0",
x"00BF",
x"00C2",
x"00C2",
x"00C0",
x"00C0",
x"00C3",
x"00C2",
x"00C4",
x"00C1",
x"0031",
x"0013",
x"0016",
x"0014",
x"0014",
x"0012",
x"0010",
x"000E",
x"000D",
x"000D",
x"000B",
x"000A",
x"000A",
x"000C",
x"000D",
x"000B",
x"000C",
x"000D",
x"000D",
x"000B",
x"000B",
x"000A",
x"000A",
x"0012",
x"0014",
x"0010",
x"0011",
x"0010",
x"000A",
x"000A",
x"000B",
x"000E",
x"000E",
x"000D",
x"0007",
x"0009",
x"000F",
x"0011",
x"0011",
x"0010",
x"0010",
x"000E",
x"0014",
x"000E",
x"0011",
x"0010",
x"000E",
x"0010",
x"0011",
x"000F",
x"000F",
x"000D",
x"000E",
x"000F",
x"0010",
x"000F",
x"000E",
x"000E",
x"000D",
x"000B",
x"000C",
x"000B",
x"000A",
x"0009",
x"0008",
x"0007",
x"0007",
x"0007",
x"0006",
x"0006",
x"0006",
x"0005",
x"0006",
x"0005",
x"0006",
x"0007",
x"0009",
x"0008",
x"0009",
x"0014",
x"0024",
x"0023",
x"0018",
x"0019",
x"0023",
x"002A",
x"0021",
x"0015",
x"0018",
x"0046",
x"0056",
x"002B",
x"003B",
x"0057",
x"0052",
x"0000",
x"0000",
x"0000",
x"0000",
x"00C0",
x"00C0",
x"00BF",
x"00C0",
x"00BD",
x"00BC",
x"00BE",
x"00BF",
x"00BE",
x"00BF",
x"00BF",
x"00BB",
x"00BC",
x"00BD",
x"00BC",
x"00BE",
x"00BE",
x"00BE",
x"00BE",
x"00C0",
x"00C0",
x"00BF",
x"00BF",
x"00BF",
x"00BF",
x"00C2",
x"00C1",
x"00C0",
x"00C1",
x"00C2",
x"00C0",
x"00C4",
x"00C1",
x"0032",
x"0014",
x"0017",
x"0015",
x"0014",
x"0011",
x"0011",
x"000E",
x"000B",
x"000C",
x"000B",
x"000A",
x"000C",
x"000D",
x"000E",
x"000B",
x"000C",
x"000D",
x"000C",
x"000A",
x"000A",
x"000A",
x"000A",
x"000D",
x"0013",
x"0011",
x"0012",
x"0012",
x"000C",
x"000C",
x"000A",
x"000D",
x"000E",
x"0009",
x"0007",
x"000D",
x"0010",
x"0011",
x"0012",
x"0011",
x"0011",
x"0013",
x"001C",
x"0009",
x"000D",
x"000F",
x"000D",
x"000E",
x"000D",
x"000B",
x"000A",
x"0009",
x"000A",
x"000B",
x"0009",
x"0008",
x"0008",
x"0009",
x"0008",
x"0008",
x"0008",
x"0008",
x"0008",
x"000A",
x"0009",
x"0009",
x"000A",
x"000A",
x"000A",
x"000C",
x"000C",
x"000C",
x"000B",
x"0009",
x"0007",
x"0007",
x"0008",
x"0008",
x"000D",
x"0038",
x"0040",
x"0037",
x"0032",
x"0029",
x"0020",
x"001F",
x"0020",
x"0018",
x"0011",
x"0034",
x"005D",
x"0027",
x"002F",
x"0054",
x"0053",
x"0000",
x"0000",
x"0000",
x"0000",
x"00BF",
x"00BF",
x"00BE",
x"00C0",
x"00BD",
x"00BE",
x"00BE",
x"00BE",
x"00BF",
x"00C0",
x"00BF",
x"00BC",
x"00BE",
x"00BE",
x"00BE",
x"00BD",
x"00BE",
x"00BF",
x"00BF",
x"00C2",
x"00C2",
x"00C1",
x"00BF",
x"00C0",
x"00C0",
x"00C0",
x"00C2",
x"00BF",
x"00C1",
x"00C2",
x"00C1",
x"00C2",
x"00C2",
x"003B",
x"0012",
x"0016",
x"0015",
x"0014",
x"0013",
x"0012",
x"000E",
x"000D",
x"000E",
x"000E",
x"000B",
x"000C",
x"000C",
x"000E",
x"000C",
x"000A",
x"000C",
x"000C",
x"000A",
x"000A",
x"000A",
x"000A",
x"000A",
x"0011",
x"0015",
x"0014",
x"0012",
x"0010",
x"000D",
x"000C",
x"000C",
x"0008",
x"0006",
x"0008",
x"000D",
x"000D",
x"000F",
x"0010",
x"000E",
x"000E",
x"000D",
x"000E",
x"000B",
x"0009",
x"000B",
x"0009",
x"000A",
x"000A",
x"0009",
x"0009",
x"000A",
x"000B",
x"000C",
x"000D",
x"000E",
x"000F",
x"0011",
x"0011",
x"0012",
x"0012",
x"0011",
x"0012",
x"0014",
x"0013",
x"0011",
x"0013",
x"0014",
x"0014",
x"0013",
x"0013",
x"0013",
x"0013",
x"0014",
x"000A",
x"0006",
x"0008",
x"0007",
x"0014",
x"0046",
x"004E",
x"0049",
x"0043",
x"0047",
x"003B",
x"0028",
x"001A",
x"0016",
x"0012",
x"0018",
x"0041",
x"0023",
x"000E",
x"001A",
x"001D",
x"0000",
x"0000",
x"0000",
x"0000",
x"00C0",
x"00C0",
x"00BF",
x"00C1",
x"00BF",
x"00BD",
x"00BF",
x"00BF",
x"00BF",
x"00C0",
x"00BF",
x"00BE",
x"00BE",
x"00BE",
x"00BD",
x"00BE",
x"00C0",
x"00C1",
x"00BF",
x"00C2",
x"00C1",
x"00BF",
x"00C1",
x"00C0",
x"00BF",
x"00C1",
x"00C2",
x"00BF",
x"00C2",
x"00C3",
x"00C1",
x"00C4",
x"00C5",
x"0042",
x"0010",
x"0013",
x"0015",
x"0014",
x"0011",
x"0010",
x"000E",
x"000D",
x"000D",
x"000C",
x"000B",
x"000C",
x"000B",
x"000D",
x"000B",
x"000A",
x"000C",
x"000C",
x"000C",
x"000D",
x"000B",
x"000C",
x"000C",
x"000C",
x"0013",
x"0016",
x"0013",
x"0011",
x"000F",
x"000E",
x"000C",
x"0009",
x"0005",
x"0008",
x"000B",
x"000B",
x"000C",
x"000C",
x"000E",
x"000E",
x"000F",
x"0011",
x"0012",
x"000D",
x"000F",
x"0009",
x"0012",
x"0011",
x"0011",
x"0012",
x"0011",
x"000F",
x"0010",
x"0011",
x"0011",
x"0010",
x"0012",
x"0011",
x"0011",
x"0013",
x"0012",
x"0011",
x"0012",
x"0012",
x"0012",
x"0014",
x"0013",
x"0013",
x"0013",
x"0011",
x"0012",
x"0014",
x"0014",
x"000A",
x"0007",
x"0009",
x"0009",
x"0026",
x"0049",
x"004B",
x"004B",
x"0046",
x"0049",
x"004E",
x"004A",
x"003F",
x"002D",
x"0022",
x"0015",
x"000F",
x"0010",
x"0015",
x"0024",
x"003E",
x"0000",
x"0000",
x"0000",
x"0000",
x"00C1",
x"00C1",
x"00C0",
x"00C0",
x"00BF",
x"00BD",
x"00BE",
x"00BF",
x"00C0",
x"00BF",
x"00BF",
x"00BE",
x"00BE",
x"00BF",
x"00BD",
x"00BF",
x"00C1",
x"00C0",
x"00C0",
x"00C2",
x"00C2",
x"00C0",
x"00C1",
x"00C0",
x"00BE",
x"00C1",
x"00C3",
x"00C0",
x"00C0",
x"00C1",
x"00C1",
x"00C5",
x"00C1",
x"0032",
x"0011",
x"0013",
x"0013",
x"0014",
x"0013",
x"0010",
x"000E",
x"000E",
x"000E",
x"000D",
x"000A",
x"000B",
x"000B",
x"000D",
x"000C",
x"000B",
x"000B",
x"000D",
x"000C",
x"000C",
x"000C",
x"000B",
x"000D",
x"000A",
x"000E",
x"0017",
x"0014",
x"0018",
x"001F",
x"001E",
x"0017",
x"000B",
x"0006",
x"0013",
x"0014",
x"0012",
x"0013",
x"0013",
x"0014",
x"0013",
x"0012",
x"0013",
x"0012",
x"0015",
x"0015",
x"0007",
x"0011",
x"0011",
x"000F",
x"0010",
x"000F",
x"0010",
x"0011",
x"000F",
x"000E",
x"000F",
x"0010",
x"000F",
x"0011",
x"0012",
x"0012",
x"0011",
x"0012",
x"0011",
x"0010",
x"0013",
x"0011",
x"0012",
x"0013",
x"0012",
x"0013",
x"0012",
x"0015",
x"000A",
x"0007",
x"0007",
x"0016",
x"0035",
x"0041",
x"003F",
x"004C",
x"004D",
x"0064",
x"007A",
x"0089",
x"0094",
x"008F",
x"0079",
x"006E",
x"006B",
x"006F",
x"008C",
x"0083",
x"0079",
x"0000",
x"0000",
x"0000",
x"0000",
x"00C2",
x"00C1",
x"00C1",
x"00C3",
x"00BF",
x"00BC",
x"00BF",
x"00C0",
x"00C1",
x"00C1",
x"00C0",
x"00BF",
x"00C0",
x"00C1",
x"00BF",
x"00BF",
x"00C2",
x"00BF",
x"00BF",
x"00C3",
x"00C2",
x"00C1",
x"00C2",
x"00C3",
x"00C2",
x"00C1",
x"00C2",
x"00C2",
x"00C4",
x"00C3",
x"00C2",
x"00C6",
x"00C2",
x"0030",
x"0011",
x"0012",
x"0013",
x"0014",
x"0013",
x"0012",
x"0012",
x"0010",
x"0012",
x"0011",
x"000E",
x"000E",
x"000D",
x"000F",
x"000F",
x"000E",
x"000D",
x"000F",
x"000B",
x"0010",
x"0012",
x"0007",
x"0009",
x"0008",
x"001E",
x"0033",
x"0033",
x"003A",
x"0031",
x"0025",
x"001C",
x"0011",
x"000B",
x"0008",
x"0009",
x"0013",
x"0015",
x"0014",
x"0013",
x"0013",
x"0011",
x"0010",
x"0010",
x"0012",
x"000F",
x"000C",
x"0012",
x"0011",
x"000F",
x"000F",
x"000F",
x"0011",
x"0011",
x"000F",
x"000D",
x"000F",
x"0010",
x"0010",
x"0011",
x"0011",
x"0012",
x"0011",
x"0011",
x"0011",
x"0012",
x"0012",
x"0012",
x"0013",
x"0013",
x"0012",
x"0012",
x"0012",
x"0012",
x"000D",
x"0010",
x"001D",
x"002E",
x"0042",
x"0060",
x"0070",
x"007F",
x"0093",
x"00A0",
x"00A0",
x"0092",
x"008D",
x"0095",
x"0094",
x"008E",
x"0092",
x"008D",
x"0087",
x"007D",
x"007F",
x"0000",
x"0000",
x"0000",
x"0000",
x"00C3",
x"00C2",
x"00BF",
x"00C3",
x"00C1",
x"00BE",
x"00C0",
x"00C1",
x"00C2",
x"00C2",
x"00C1",
x"00BF",
x"00C0",
x"00C0",
x"00C0",
x"00C0",
x"00C2",
x"00C0",
x"00C2",
x"00C3",
x"00C2",
x"00C3",
x"00C3",
x"00C1",
x"00C1",
x"00C3",
x"00C4",
x"00C3",
x"00C4",
x"00C5",
x"00C2",
x"00C6",
x"00C0",
x"002E",
x"0010",
x"0012",
x"0013",
x"0013",
x"0012",
x"0011",
x"0011",
x"0011",
x"0012",
x"0011",
x"000E",
x"000F",
x"000F",
x"0010",
x"0011",
x"0010",
x"000E",
x"000C",
x"000A",
x"000F",
x"000C",
x"0009",
x"0006",
x"0008",
x"0022",
x"003A",
x"0038",
x"0039",
x"002D",
x"0020",
x"0023",
x"0019",
x"0010",
x"0008",
x"0008",
x"0010",
x"0014",
x"0013",
x"0011",
x"0012",
x"0012",
x"0013",
x"000F",
x"000F",
x"000C",
x"000C",
x"0010",
x"000F",
x"0010",
x"0012",
x"0011",
x"0010",
x"0011",
x"000F",
x"000E",
x"000F",
x"0011",
x"000F",
x"000E",
x"0011",
x"0010",
x"0011",
x"0010",
x"0010",
x"0010",
x"0010",
x"0010",
x"000E",
x"000F",
x"000E",
x"0009",
x"0010",
x"0019",
x"0052",
x"007D",
x"0078",
x"007A",
x"0088",
x"0097",
x"009F",
x"00A0",
x"0097",
x"009C",
x"0098",
x"0086",
x"008A",
x"008F",
x"008E",
x"0089",
x"0085",
x"008A",
x"0086",
x"008D",
x"008B",
x"0000",
x"0000",
x"0000",
x"0000",
x"00C3",
x"00C3",
x"00C1",
x"00C3",
x"00C2",
x"00C0",
x"00C1",
x"00C2",
x"00C0",
x"00C2",
x"00C1",
x"00C0",
x"00C1",
x"00C2",
x"00C0",
x"00C0",
x"00C1",
x"00BF",
x"00C1",
x"00C4",
x"00C3",
x"00C1",
x"00C3",
x"00C3",
x"00C1",
x"00C3",
x"00C5",
x"00C4",
x"00C5",
x"00C5",
x"00C4",
x"00CA",
x"00B9",
x"0022",
x"0010",
x"0011",
x"0011",
x"0012",
x"0011",
x"0012",
x"0012",
x"0011",
x"0010",
x"0013",
x"000E",
x"000F",
x"0010",
x"0011",
x"000F",
x"000F",
x"000F",
x"000C",
x"000A",
x"0009",
x"0009",
x"000D",
x"000A",
x"0020",
x"001C",
x"0035",
x"003A",
x"003D",
x"0031",
x"002B",
x"002B",
x"0020",
x"0016",
x"0011",
x"0007",
x"000C",
x"0012",
x"0013",
x"0012",
x"0011",
x"0011",
x"000F",
x"000F",
x"000E",
x"0011",
x"0009",
x"0010",
x"000F",
x"000E",
x"0011",
x"0011",
x"0010",
x"000F",
x"0010",
x"0010",
x"0011",
x"0011",
x"000F",
x"000F",
x"0011",
x"0010",
x"0011",
x"0010",
x"0010",
x"000C",
x"000C",
x"000A",
x"000F",
x"001D",
x"0031",
x"004F",
x"0069",
x"0082",
x"0082",
x"0090",
x"008A",
x"0088",
x"0090",
x"0093",
x"0096",
x"0097",
x"008B",
x"009C",
x"009E",
x"0089",
x"0088",
x"008B",
x"008D",
x"008B",
x"0085",
x"008A",
x"008E",
x"009D",
x"008A",
x"0000",
x"0000",
x"0000",
x"0000",
x"00C2",
x"00C2",
x"00C3",
x"00C4",
x"00C0",
x"00C0",
x"00C2",
x"00C2",
x"00C0",
x"00C2",
x"00C2",
x"00C2",
x"00C2",
x"00C2",
x"00BF",
x"00C0",
x"00C1",
x"00C1",
x"00C2",
x"00C5",
x"00C2",
x"00C2",
x"00C4",
x"00C4",
x"00C0",
x"00C3",
x"00C4",
x"00C4",
x"00C5",
x"00C5",
x"00C6",
x"00D1",
x"00A5",
x"0018",
x"0010",
x"0010",
x"0010",
x"0013",
x"0012",
x"0011",
x"0011",
x"0011",
x"0013",
x"0033",
x"0014",
x"000A",
x"000E",
x"0010",
x"000B",
x"0008",
x"000E",
x"000C",
x"000A",
x"0009",
x"0008",
x"0007",
x"0038",
x"0043",
x"0008",
x"001E",
x"0045",
x"004A",
x"003B",
x"0033",
x"002B",
x"0025",
x"0019",
x"0029",
x"000E",
x"0006",
x"000F",
x"0011",
x"000F",
x"000E",
x"0010",
x"000E",
x"000D",
x"000F",
x"0012",
x"000B",
x"000F",
x"000F",
x"000D",
x"0010",
x"0011",
x"000F",
x"0010",
x"0011",
x"000F",
x"0010",
x"000F",
x"000F",
x"000E",
x"0010",
x"000C",
x"000B",
x"000B",
x"000D",
x"001B",
x"002F",
x"0045",
x"006C",
x"0094",
x"00A1",
x"00AD",
x"00A6",
x"0092",
x"0083",
x"0091",
x"0085",
x"007B",
x"0082",
x"0089",
x"0091",
x"00A1",
x"0096",
x"00A0",
x"0093",
x"008E",
x"0095",
x"0092",
x"0090",
x"0087",
x"0093",
x"008A",
x"0086",
x"0080",
x"0096",
x"0000",
x"0000",
x"0000",
x"0000",
x"00C2",
x"00C1",
x"00C3",
x"00C4",
x"00BF",
x"00C0",
x"00C2",
x"00C0",
x"00C0",
x"00C3",
x"00C3",
x"00C1",
x"00C1",
x"00C1",
x"00BE",
x"00BF",
x"00C3",
x"00C2",
x"00C2",
x"00C4",
x"00C3",
x"00C2",
x"00C3",
x"00C4",
x"00C1",
x"00C4",
x"00C5",
x"00C5",
x"00CC",
x"00CF",
x"00CC",
x"00B6",
x"0042",
x"0009",
x"000E",
x"000D",
x"000D",
x"0013",
x"0016",
x"000A",
x"000A",
x"0011",
x"0011",
x"001F",
x"001B",
x"000D",
x"000D",
x"0012",
x"000B",
x"0007",
x"000C",
x"000C",
x"000A",
x"000B",
x"0009",
x"000A",
x"004A",
x"0021",
x"000F",
x"000C",
x"0039",
x"0048",
x"0032",
x"002A",
x"0028",
x"002A",
x"0015",
x"0018",
x"0021",
x"0008",
x"000D",
x"0010",
x"000F",
x"0010",
x"000F",
x"0011",
x"0010",
x"0011",
x"0011",
x"000D",
x"0011",
x"0012",
x"000F",
x"0011",
x"0011",
x"0010",
x"0011",
x"000F",
x"000D",
x"0010",
x"000F",
x"0010",
x"000C",
x"0008",
x"0019",
x"002B",
x"0049",
x"005C",
x"008D",
x"00A5",
x"009C",
x"00A6",
x"00A0",
x"009F",
x"0098",
x"0097",
x"0093",
x"0080",
x"0098",
x"0083",
x"0071",
x"008C",
x"008B",
x"008D",
x"0096",
x"008A",
x"009B",
x"008B",
x"0085",
x"008D",
x"009E",
x"0083",
x"0080",
x"0094",
x"0095",
x"0094",
x"0087",
x"008A",
x"0000",
x"0000",
x"0000",
x"0000",
x"00C4",
x"00C3",
x"00C1",
x"00C4",
x"00C0",
x"00C0",
x"00C1",
x"00C1",
x"00C1",
x"00C3",
x"00C4",
x"00C3",
x"00C3",
x"00C0",
x"00BF",
x"00BF",
x"00C3",
x"00C2",
x"00C2",
x"00C5",
x"00C5",
x"00C2",
x"00C4",
x"00C5",
x"00C6",
x"00C9",
x"00CF",
x"00C7",
x"009D",
x"0095",
x"0065",
x"0023",
x"0004",
x"0006",
x"0005",
x"0006",
x"0007",
x"0008",
x"0007",
x"0007",
x"0008",
x"0010",
x"0011",
x"000E",
x"000F",
x"0012",
x"0013",
x"0011",
x"000C",
x"0008",
x"000A",
x"000B",
x"000C",
x"000C",
x"0009",
x"0009",
x"000F",
x"000F",
x"000E",
x"0007",
x"0024",
x"0039",
x"0019",
x"0024",
x"0020",
x"001E",
x"0022",
x"000B",
x"001F",
x"0013",
x"000D",
x"0011",
x"0013",
x"0011",
x"0012",
x"0010",
x"000F",
x"000F",
x"0010",
x"000B",
x"000E",
x"0010",
x"000E",
x"0010",
x"000F",
x"0010",
x"0010",
x"000F",
x"000B",
x"000A",
x"000A",
x"0007",
x"0024",
x"0058",
x"0087",
x"008D",
x"009B",
x"0098",
x"009F",
x"00A3",
x"0092",
x"009A",
x"009D",
x"0098",
x"0094",
x"0094",
x"008E",
x"0083",
x"008E",
x"007E",
x"007C",
x"0088",
x"008E",
x"0098",
x"0097",
x"0092",
x"0096",
x"008B",
x"008F",
x"0097",
x"009A",
x"0080",
x"007D",
x"0087",
x"009B",
x"008B",
x"0093",
x"008A",
x"0000",
x"0000",
x"0000",
x"0000",
x"00C2",
x"00C2",
x"00C1",
x"00C3",
x"00C0",
x"00C0",
x"00C2",
x"00C2",
x"00C1",
x"00C4",
x"00C4",
x"00C2",
x"00C2",
x"00C1",
x"00C1",
x"00C0",
x"00C3",
x"00C4",
x"00C2",
x"00C5",
x"00C7",
x"00C6",
x"00CA",
x"00CF",
x"00C3",
x"00B1",
x"00A1",
x"0068",
x"000F",
x"0010",
x"0008",
x"000A",
x"000C",
x"000D",
x"0010",
x"0006",
x"0000",
x"0000",
x"0003",
x"0005",
x"0006",
x"000A",
x"000C",
x"0007",
x"0006",
x"0008",
x"0009",
x"000B",
x"000B",
x"0009",
x"000B",
x"000A",
x"000A",
x"000B",
x"0001",
x"0036",
x"0049",
x"000C",
x"000A",
x"0009",
x"001D",
x"0023",
x"000B",
x"001B",
x"0026",
x"000E",
x"0021",
x"000D",
x"000B",
x"0012",
x"0012",
x"0012",
x"0012",
x"0011",
x"0012",
x"0010",
x"000F",
x"0010",
x"000C",
x"0007",
x"000C",
x"000E",
x"000D",
x"000E",
x"000B",
x"0008",
x"0004",
x"000A",
x"0017",
x"0022",
x"0030",
x"0051",
x"0089",
x"00A5",
x"009E",
x"008E",
x"0096",
x"0094",
x"009E",
x"00A3",
x"0094",
x"009B",
x"00A4",
x"009B",
x"009A",
x"0099",
x"008E",
x"007F",
x"0087",
x"0069",
x"0093",
x"0088",
x"008E",
x"0092",
x"008F",
x"0091",
x"0096",
x"0094",
x"009B",
x"00A0",
x"00A5",
x"0088",
x"007B",
x"0076",
x"0069",
x"0059",
x"0048",
x"003C",
x"0000",
x"0000",
x"0000",
x"0000",
x"00C1",
x"00C1",
x"00C3",
x"00C5",
x"00C1",
x"00C1",
x"00C4",
x"00C2",
x"00C2",
x"00C4",
x"00C4",
x"00C3",
x"00C3",
x"00C3",
x"00C2",
x"00C1",
x"00C4",
x"00C4",
x"00C4",
x"00C7",
x"00C7",
x"00C3",
x"00C6",
x"007B",
x"003B",
x"001C",
x"0011",
x"000B",
x"0004",
x"0006",
x"0008",
x"0008",
x"0009",
x"000F",
x"0047",
x"007B",
x"0070",
x"004E",
x"001E",
x"0006",
x"0005",
x"0015",
x"0015",
x"000A",
x"0007",
x"0006",
x"0006",
x"0008",
x"000A",
x"000B",
x"000A",
x"000A",
x"000A",
x"0003",
x"0041",
x"008D",
x"0039",
x"000C",
x"000D",
x"000A",
x"000D",
x"000C",
x"000D",
x"0010",
x"001B",
x"000E",
x"001A",
x"0028",
x"0013",
x"000A",
x"0010",
x"0012",
x"0011",
x"0012",
x"0011",
x"0010",
x"000F",
x"000F",
x"000A",
x"0008",
x"000B",
x"000B",
x"0009",
x"0006",
x"0010",
x"002E",
x"0071",
x"0077",
x"0071",
x"0097",
x"0094",
x"00AB",
x"00A2",
x"0095",
x"0096",
x"0091",
x"0098",
x"0096",
x"009D",
x"00A7",
x"0099",
x"009F",
x"00A1",
x"009D",
x"00A3",
x"00A2",
x"0093",
x"0080",
x"008B",
x"006F",
x"008A",
x"0089",
x"008E",
x"0093",
x"0091",
x"0090",
x"009A",
x"0098",
x"0086",
x"0076",
x"0066",
x"004A",
x"003A",
x"0031",
x"0031",
x"003D",
x"004A",
x"005B",
x"0000",
x"0000",
x"0000",
x"0000",
x"00C3",
x"00C2",
x"00C3",
x"00C5",
x"00C2",
x"00C1",
x"00C4",
x"00C3",
x"00C2",
x"00C3",
x"00C5",
x"00C2",
x"00C4",
x"00C4",
x"00C2",
x"00C3",
x"00C4",
x"00C5",
x"00C5",
x"00D2",
x"0093",
x"004D",
x"0046",
x"000A",
x"0003",
x"0004",
x"0007",
x"0008",
x"0007",
x"0007",
x"0008",
x"0007",
x"0006",
x"0026",
x"004E",
x"007A",
x"00C3",
x"00DF",
x"00AC",
x"005E",
x"0055",
x"0021",
x"0012",
x"000C",
x"0007",
x"0009",
x"000E",
x"000B",
x"0010",
x"000A",
x"0009",
x"000A",
x"0005",
x"004E",
x"008B",
x"002B",
x"0003",
x"0012",
x"000F",
x"000B",
x"000A",
x"000A",
x"000D",
x"000E",
x"0011",
x"0011",
x"0014",
x"0031",
x"001B",
x"000D",
x"000E",
x"0011",
x"0011",
x"0012",
x"0011",
x"0010",
x"000E",
x"000F",
x"000D",
x"000E",
x"000A",
x"0009",
x"0010",
x"003D",
x"0082",
x"00A5",
x"00F4",
x"00C1",
x"0087",
x"00A3",
x"0099",
x"00A7",
x"009B",
x"0097",
x"0096",
x"0092",
x"0095",
x"0092",
x"009E",
x"00AB",
x"0092",
x"009B",
x"00A2",
x"0099",
x"00A6",
x"00A7",
x"0099",
x"007B",
x"0091",
x"0086",
x"008C",
x"007E",
x"0079",
x"0066",
x"005E",
x"0064",
x"0056",
x"0044",
x"0037",
x"0032",
x"0036",
x"0047",
x"005C",
x"0072",
x"0088",
x"00A5",
x"00BD",
x"00C9",
x"0000",
x"0000",
x"0000",
x"0000",
x"00C4",
x"00C4",
x"00C4",
x"00C6",
x"00C3",
x"00C2",
x"00C4",
x"00C3",
x"00C3",
x"00C6",
x"00C3",
x"00C4",
x"00C4",
x"00C4",
x"00C3",
x"00C4",
x"00C3",
x"00C6",
x"00CC",
x"00B5",
x"0025",
x"0006",
x"0005",
x"0008",
x"0008",
x"0007",
x"000A",
x"000A",
x"0008",
x"0007",
x"0007",
x"0008",
x"000A",
x"003E",
x"0066",
x"006A",
x"0080",
x"00B7",
x"00B5",
x"0085",
x"009E",
x"0084",
x"0079",
x"006A",
x"005C",
x"006A",
x"0027",
x"0016",
x"000E",
x"0007",
x"000A",
x"0006",
x"0056",
x"0087",
x"001E",
x"0006",
x"0009",
x"0011",
x"000E",
x"000A",
x"000A",
x"000C",
x"000D",
x"000F",
x"0012",
x"0013",
x"0011",
x"0015",
x"0013",
x"000F",
x"0010",
x"0010",
x"000F",
x"000F",
x"000F",
x"000D",
x"0006",
x"000B",
x"0018",
x"001B",
x"002F",
x"004A",
x"001B",
x"006B",
x"00B3",
x"00A9",
x"00EF",
x"00B3",
x"0083",
x"00A2",
x"0098",
x"00A9",
x"009C",
x"0099",
x"0097",
x"0090",
x"0096",
x"0097",
x"009E",
x"00A5",
x"008B",
x"0094",
x"00A3",
x"009F",
x"00A6",
x"00AB",
x"009C",
x"007F",
x"0071",
x"0054",
x"003F",
x"0022",
x"0030",
x"004F",
x"0044",
x"0048",
x"006B",
x"0056",
x"0070",
x"0089",
x"00A0",
x"00B6",
x"00CC",
x"00E0",
x"00ED",
x"00F6",
x"00FC",
x"00F9",
x"0000",
x"0000",
x"0000",
x"0000",
x"00C5",
x"00C5",
x"00C5",
x"00C8",
x"00C3",
x"00C3",
x"00C5",
x"00C4",
x"00C3",
x"00C6",
x"00C5",
x"00C4",
x"00C4",
x"00C5",
x"00C3",
x"00C3",
x"00C4",
x"00C7",
x"00CB",
x"0071",
x"000B",
x"000F",
x"0009",
x"0008",
x"0008",
x"0008",
x"0008",
x"0008",
x"0005",
x"0004",
x"0007",
x"000B",
x"0013",
x"0023",
x"0052",
x"008B",
x"0086",
x"0082",
x"00AD",
x"00B1",
x"0089",
x"006E",
x"006E",
x"0053",
x"0060",
x"003B",
x"001C",
x"0016",
x"0009",
x"000C",
x"0006",
x"0055",
x"0079",
x"0018",
x"0004",
x"000B",
x"000C",
x"0012",
x"000B",
x"0008",
x"000A",
x"000D",
x"000F",
x"0011",
x"0013",
x"0012",
x"0011",
x"000E",
x"000C",
x"000D",
x"000E",
x"000F",
x"000C",
x"000A",
x"0008",
x"0016",
x"0055",
x"008D",
x"00BB",
x"00AD",
x"00A7",
x"0094",
x"0022",
x"0070",
x"00B1",
x"00AD",
x"00EF",
x"00BA",
x"008F",
x"00A1",
x"0099",
x"00A9",
x"009E",
x"009C",
x"0099",
x"0090",
x"009B",
x"009C",
x"00A0",
x"00AA",
x"0090",
x"009A",
x"0096",
x"0086",
x"006F",
x"0057",
x"0034",
x"0018",
x"000F",
x"0004",
x"0003",
x"0000",
x"001B",
x"002F",
x"0090",
x"00DB",
x"00EE",
x"00C8",
x"00DC",
x"00EE",
x"00F6",
x"00F8",
x"00F7",
x"00F1",
x"00DD",
x"00C1",
x"00B0",
x"0098",
x"0000",
x"0000",
x"0000",
x"0000",
x"00C5",
x"00C5",
x"00C7",
x"00C7",
x"00C4",
x"00C4",
x"00C5",
x"00C3",
x"00C3",
x"00C6",
x"00C6",
x"00C3",
x"00C5",
x"00C7",
x"00C3",
x"00C4",
x"00C5",
x"00CA",
x"00BE",
x"0035",
x"0010",
x"000D",
x"0007",
x"0006",
x"0007",
x"0008",
x"0008",
x"0005",
x"001B",
x"006D",
x"0074",
x"0060",
x"002E",
x"0016",
x"0021",
x"005A",
x"0074",
x"0067",
x"0093",
x"00A0",
x"0067",
x"004C",
x"0021",
x"000B",
x"0013",
x"0017",
x"001C",
x"000F",
x"000A",
x"000E",
x"0064",
x"0069",
x"0014",
x"000D",
x"0009",
x"0008",
x"000D",
x"000E",
x"0009",
x"000A",
x"000A",
x"000F",
x"0013",
x"0013",
x"0013",
x"0010",
x"000E",
x"000D",
x"000C",
x"000C",
x"000A",
x"0005",
x"000D",
x"002A",
x"006B",
x"00A0",
x"00C9",
x"00DA",
x"00E2",
x"00C2",
x"00AE",
x"008E",
x"0024",
x"0067",
x"00A6",
x"00AD",
x"00F0",
x"00BC",
x"0096",
x"00A1",
x"009C",
x"00AA",
x"00A0",
x"009E",
x"009E",
x"0096",
x"00A3",
x"00A4",
x"00A0",
x"0084",
x"004D",
x"003B",
x"002A",
x"001E",
x"000A",
x"0002",
x"0001",
x"0002",
x"0002",
x"0003",
x"0009",
x"001A",
x"0026",
x"0049",
x"00C5",
x"00EE",
x"00FE",
x"00EE",
x"00EB",
x"00D7",
x"00BE",
x"00A9",
x"0096",
x"0086",
x"0090",
x"0092",
x"0086",
x"0085",
x"0000",
x"0000",
x"0000",
x"0000",
x"00C3",
x"00C3",
x"00C5",
x"00C5",
x"00C3",
x"00C3",
x"00C5",
x"00C4",
x"00C3",
x"00C6",
x"00C6",
x"00C5",
x"00C6",
x"00C5",
x"00C4",
x"00C5",
x"00C6",
x"00CE",
x"00A2",
x"0010",
x"000B",
x"000B",
x"0007",
x"0006",
x"0007",
x"0007",
x"0006",
x"000A",
x"0050",
x"009A",
x"0087",
x"0086",
x"00A6",
x"0043",
x"001D",
x"003F",
x"0045",
x"0044",
x"006F",
x"008E",
x"0066",
x"004A",
x"0010",
x"0013",
x"0014",
x"001A",
x"0014",
x"0006",
x"000D",
x"0077",
x"006D",
x"0011",
x"000D",
x"0011",
x"0009",
x"000B",
x"000D",
x"000B",
x"000B",
x"000B",
x"000D",
x"0012",
x"0013",
x"0011",
x"0010",
x"000D",
x"000A",
x"000A",
x"0006",
x"0008",
x"0020",
x"0059",
x"008E",
x"00AB",
x"00B7",
x"00B5",
x"00C8",
x"00D0",
x"00DD",
x"00BD",
x"00A9",
x"0084",
x"0020",
x"0068",
x"0096",
x"00B2",
x"00F3",
x"00B5",
x"0091",
x"00A3",
x"00A6",
x"00B6",
x"00A9",
x"00A2",
x"008F",
x"0068",
x"0051",
x"0037",
x"001E",
x"0010",
x"0004",
x"0000",
x"003F",
x"0052",
x"0005",
x"000A",
x"001C",
x"0034",
x"005B",
x"007F",
x"008C",
x"008A",
x"006E",
x"0052",
x"0085",
x"00E9",
x"00F6",
x"00C0",
x"008E",
x"009E",
x"0094",
x"0076",
x"007B",
x"0081",
x"009B",
x"0097",
x"0092",
x"0085",
x"0000",
x"0000",
x"0000",
x"0000",
x"00C5",
x"00C4",
x"00C5",
x"00C6",
x"00C1",
x"00C3",
x"00C5",
x"00C3",
x"00C3",
x"00C7",
x"00C5",
x"00C6",
x"00C6",
x"00C6",
x"00C4",
x"00C5",
x"00C7",
x"00D1",
x"008A",
x"0002",
x"000A",
x"000B",
x"0008",
x"0008",
x"0008",
x"0007",
x"0007",
x"000C",
x"0036",
x"0035",
x"007E",
x"0074",
x"0095",
x"0077",
x"0037",
x"0017",
x"0015",
x"0019",
x"0029",
x"0043",
x"0034",
x"0018",
x"000C",
x"0016",
x"0014",
x"0019",
x"000C",
x"000C",
x"0074",
x"0076",
x"0011",
x"000E",
x"0010",
x"000D",
x"000B",
x"000B",
x"000A",
x"000E",
x"0010",
x"000B",
x"0010",
x"0013",
x"0012",
x"000D",
x"000D",
x"0009",
x"0006",
x"0012",
x"003F",
x"007A",
x"00A8",
x"00BB",
x"00BA",
x"00B5",
x"00BB",
x"00AD",
x"00C5",
x"00D1",
x"00DD",
x"00BB",
x"00A9",
x"0085",
x"001C",
x"0067",
x"0093",
x"00A7",
x"00FA",
x"00C1",
x"0098",
x"00A1",
x"008F",
x"0072",
x"0051",
x"002C",
x"0013",
x"0008",
x"0001",
x"0000",
x"0000",
x"0002",
x"0009",
x"0016",
x"0099",
x"00C6",
x"007E",
x"008A",
x"0088",
x"007D",
x"0067",
x"0045",
x"0032",
x"002D",
x"0041",
x"0050",
x"0066",
x"00A1",
x"009E",
x"00A3",
x"0095",
x"0095",
x"0093",
x"007D",
x"0084",
x"009A",
x"009A",
x"0085",
x"008E",
x"0085",
x"0000",
x"0000",
x"0000",
x"0000",
x"00C3",
x"00C3",
x"00C4",
x"00C8",
x"00C4",
x"00C1",
x"00C4",
x"00C2",
x"00C3",
x"00C7",
x"00C4",
x"00C4",
x"00C6",
x"00C7",
x"00C5",
x"00C5",
x"00C6",
x"00D0",
x"0092",
x"0005",
x"000A",
x"000C",
x"000D",
x"000E",
x"000A",
x"0009",
x"000A",
x"0009",
x"0009",
x"0012",
x"0084",
x"008C",
x"0080",
x"0083",
x"0071",
x"003D",
x"0014",
x"000F",
x"0012",
x"000D",
x"0006",
x"0005",
x"0008",
x"0014",
x"001A",
x"000E",
x"0014",
x"0078",
x"006A",
x"000C",
x"000E",
x"0010",
x"000D",
x"000E",
x"000C",
x"000B",
x"000D",
x"0012",
x"000E",
x"000C",
x"0011",
x"0011",
x"000E",
x"000A",
x"000C",
x"0033",
x"006E",
x"009F",
x"00B7",
x"00BD",
x"00B7",
x"00B5",
x"00B4",
x"00B7",
x"00C6",
x"00B0",
x"00C7",
x"00D3",
x"00DF",
x"00BB",
x"00AE",
x"0088",
x"0017",
x"0062",
x"00A6",
x"00A6",
x"00B6",
x"006C",
x"0036",
x"001F",
x"000E",
x"0002",
x"0000",
x"0000",
x"0002",
x"0008",
x"001A",
x"002A",
x"004B",
x"006E",
x"007C",
x"007D",
x"00B1",
x"00E9",
x"005F",
x"002F",
x"0038",
x"003E",
x"0049",
x"005B",
x"0080",
x"0080",
x"0090",
x"00A5",
x"0090",
x"0087",
x"0091",
x"0092",
x"0097",
x"0097",
x"0080",
x"007D",
x"0081",
x"008D",
x"0095",
x"0083",
x"0086",
x"0086",
x"0000",
x"0000",
x"0000",
x"0000",
x"00C3",
x"00C3",
x"00C5",
x"00C7",
x"00C3",
x"00C3",
x"00C4",
x"00C3",
x"00C3",
x"00C7",
x"00C4",
x"00C4",
x"00C6",
x"00C6",
x"00C5",
x"00C6",
x"00C8",
x"00CD",
x"00AA",
x"0011",
x"0008",
x"000B",
x"000B",
x"000F",
x"000A",
x"000A",
x"000A",
x"0008",
x"0007",
x"0006",
x"000C",
x"0010",
x"005D",
x"00A1",
x"0094",
x"0070",
x"0039",
x"0010",
x"000E",
x"000B",
x"0006",
x"0006",
x"0006",
x"000A",
x"0011",
x"0015",
x"007E",
x"005F",
x"0008",
x"0009",
x"000F",
x"000D",
x"000D",
x"000E",
x"000E",
x"000D",
x"0010",
x"0011",
x"000E",
x"0010",
x"000E",
x"000C",
x"000A",
x"0009",
x"0006",
x"0047",
x"00B7",
x"00BD",
x"00B5",
x"00B6",
x"00B4",
x"00B5",
x"00B4",
x"00B7",
x"00C8",
x"00B5",
x"00CE",
x"00DC",
x"00E7",
x"00BE",
x"00A9",
x"0078",
x"0019",
x"0031",
x"002E",
x"0016",
x"0009",
x"0000",
x"0000",
x"0001",
x"000A",
x"001A",
x"0029",
x"0049",
x"0073",
x"007E",
x"0083",
x"0079",
x"005F",
x"0038",
x"002D",
x"003C",
x"0081",
x"009C",
x"0076",
x"007C",
x"009C",
x"0077",
x"006D",
x"007C",
x"0095",
x"0085",
x"007B",
x"008F",
x"0095",
x"008F",
x"0091",
x"009B",
x"0091",
x"008A",
x"008D",
x"0082",
x"0084",
x"0093",
x"008F",
x"0090",
x"008D",
x"007A",
x"0000",
x"0000",
x"0000",
x"0000",
x"00C4",
x"00C5",
x"00C6",
x"00C7",
x"00C4",
x"00C3",
x"00C5",
x"00C3",
x"00C3",
x"00C7",
x"00C5",
x"00C4",
x"00C6",
x"00C7",
x"00C5",
x"00C7",
x"00C8",
x"00CB",
x"00BA",
x"001B",
x"0008",
x"000C",
x"000C",
x"000B",
x"000B",
x"000B",
x"000A",
x"0009",
x"0006",
x"0013",
x"003F",
x"0053",
x"0087",
x"00A8",
x"00A2",
x"008E",
x"006A",
x"0037",
x"000D",
x"000A",
x"0006",
x"0007",
x"0008",
x"0006",
x"000A",
x"0080",
x"0054",
x"000C",
x"000C",
x"000A",
x"0009",
x"000C",
x"000B",
x"000F",
x"000D",
x"000F",
x"000F",
x"000D",
x"000C",
x"000C",
x"0008",
x"0008",
x"0007",
x"0007",
x"0007",
x"0002",
x"004F",
x"00B9",
x"00B7",
x"00B5",
x"00B7",
x"00B9",
x"00BD",
x"00C8",
x"00CF",
x"00B3",
x"00B2",
x"0096",
x"0076",
x"0046",
x"001A",
x"000C",
x"0004",
x"0000",
x"0000",
x"0008",
x"001E",
x"002F",
x"0052",
x"006F",
x"0072",
x"0074",
x"0070",
x"005E",
x"0045",
x"0026",
x"0013",
x"0016",
x"0031",
x"0071",
x"00A4",
x"00B4",
x"00A6",
x"0096",
x"009B",
x"009C",
x"00A3",
x"006F",
x"005C",
x"0090",
x"0091",
x"008A",
x"007C",
x"008B",
x"008C",
x"0093",
x"0095",
x"0092",
x"008E",
x"008F",
x"00A1",
x"0085",
x"0087",
x"0097",
x"0091",
x"0094",
x"0093",
x"0073",
x"0000",
x"0000",
x"0000",
x"0000",
x"00C5",
x"00C5",
x"00C5",
x"00C6",
x"00C5",
x"00C3",
x"00C5",
x"00C5",
x"00C5",
x"00C7",
x"00C4",
x"00C4",
x"00C6",
x"00C7",
x"00C6",
x"00C6",
x"00C6",
x"00C9",
x"00C4",
x"002A",
x"0006",
x"000A",
x"000C",
x"000F",
x"000B",
x"0009",
x"0009",
x"0007",
x"000D",
x"007E",
x"00C3",
x"00BA",
x"00AD",
x"00AE",
x"00AD",
x"009A",
x"0082",
x"0062",
x"002B",
x"0007",
x"0001",
x"0003",
x"0007",
x"0004",
x"0048",
x"0079",
x"000F",
x"000E",
x"0011",
x"000E",
x"0007",
x"0009",
x"0009",
x"000C",
x"000D",
x"000C",
x"000C",
x"000A",
x"000A",
x"0007",
x"0006",
x"0006",
x"0006",
x"0006",
x"0006",
x"0004",
x"0008",
x"0077",
x"00C5",
x"00BF",
x"00B5",
x"00A9",
x"0090",
x"007B",
x"005B",
x"0025",
x"000F",
x"0005",
x"0000",
x"0000",
x"000E",
x"0021",
x"002F",
x"0045",
x"0059",
x"0063",
x"0078",
x"007A",
x"005A",
x"003B",
x"0037",
x"0041",
x"004E",
x"004C",
x"0047",
x"002E",
x"004E",
x"0089",
x"00B8",
x"00BA",
x"0097",
x"0099",
x"0098",
x"009A",
x"0094",
x"0095",
x"009D",
x"0079",
x"0076",
x"0095",
x"008E",
x"0086",
x"007F",
x"0086",
x"0094",
x"008A",
x"0087",
x"0094",
x"008C",
x"0092",
x"0098",
x"0081",
x"0080",
x"0091",
x"0081",
x"008E",
x"0095",
x"0090",
x"0000",
x"0000",
x"0000",
x"0000",
x"00C5",
x"00C5",
x"00C7",
x"00C9",
x"00C6",
x"00C5",
x"00C6",
x"00C5",
x"00C5",
x"00C6",
x"00C5",
x"00C4",
x"00C7",
x"00C9",
x"00C6",
x"00C6",
x"00C5",
x"00C6",
x"00CD",
x"0059",
x"0002",
x"000B",
x"000E",
x"000E",
x"000B",
x"0007",
x"0007",
x"0007",
x"0051",
x"00C2",
x"00B9",
x"00C8",
x"00BC",
x"00B8",
x"00BC",
x"00AB",
x"0086",
x"007A",
x"006D",
x"002F",
x"003A",
x"001E",
x"000A",
x"0004",
x"0077",
x"0042",
x"0007",
x"0010",
x"000F",
x"000F",
x"000B",
x"0007",
x"0008",
x"0006",
x"0008",
x"0008",
x"0008",
x"0007",
x"0007",
x"0006",
x"0007",
x"0006",
x"0006",
x"0006",
x"0006",
x"0006",
x"0003",
x"001B",
x"0072",
x"0063",
x"0036",
x"0014",
x"0005",
x"0000",
x"0000",
x"0014",
x"002B",
x"0031",
x"0046",
x"0057",
x"005E",
x"006E",
x"006E",
x"0055",
x"0043",
x"003C",
x"005D",
x"0064",
x"006A",
x"0086",
x"00A3",
x"009B",
x"006C",
x"0049",
x"0064",
x"00A3",
x"00BD",
x"00AE",
x"009E",
x"009B",
x"0084",
x"0090",
x"0099",
x"00A1",
x"009A",
x"0095",
x"0099",
x"007A",
x"0079",
x"0087",
x"008A",
x"0089",
x"0082",
x"008C",
x"009E",
x"008F",
x"0088",
x"0096",
x"0094",
x"0096",
x"008C",
x"0083",
x"007D",
x"0093",
x"008D",
x"0091",
x"0096",
x"0078",
x"0000",
x"0000",
x"0000",
x"0000",
x"00C5",
x"00C5",
x"00C7",
x"00C9",
x"00C6",
x"00C7",
x"00C7",
x"00C5",
x"00C6",
x"00C7",
x"00C6",
x"00C3",
x"00C6",
x"00C9",
x"00C7",
x"00C7",
x"00C6",
x"00C4",
x"00CE",
x"00A4",
x"0013",
x"0007",
x"000C",
x"000D",
x"000B",
x"0006",
x"0005",
x"0018",
x"009B",
x"00B8",
x"007C",
x"00B7",
x"00BE",
x"00BE",
x"00B1",
x"0092",
x"007E",
x"0089",
x"0083",
x"0070",
x"00C0",
x"00BB",
x"007D",
x"0025",
x"0082",
x"0031",
x"000D",
x"0006",
x"0008",
x"0008",
x"0008",
x"0008",
x"0008",
x"0006",
x"0007",
x"0006",
x"0006",
x"0007",
x"0008",
x"0006",
x"0006",
x"0006",
x"0006",
x"0007",
x"0008",
x"0006",
x"0004",
x"0002",
x"0000",
x"0000",
x"0015",
x"0026",
x"0033",
x"004B",
x"004F",
x"005A",
x"0076",
x"0062",
x"0042",
x"0038",
x"003E",
x"0031",
x"002D",
x"0073",
x"009B",
x"008A",
x"0093",
x"0096",
x"00A4",
x"0090",
x"006D",
x"0052",
x"0073",
x"00AD",
x"00BF",
x"00A3",
x"0090",
x"008B",
x"009F",
x"009A",
x"0080",
x"009A",
x"009B",
x"00A1",
x"00A2",
x"009B",
x"0094",
x"007A",
x"0083",
x"0086",
x"0086",
x"009A",
x"0095",
x"009D",
x"009B",
x"0091",
x"008B",
x"0097",
x"009F",
x"00A2",
x"009D",
x"0089",
x"007F",
x"0090",
x"0099",
x"0096",
x"0097",
x"0085",
x"0000",
x"0000",
x"0000",
x"0000",
x"00C4",
x"00C5",
x"00C7",
x"00C9",
x"00C6",
x"00C4",
x"00C6",
x"00C5",
x"00C5",
x"00C7",
x"00C5",
x"00C4",
x"00C7",
x"00C8",
x"00C6",
x"00C6",
x"00C5",
x"00C4",
x"00CA",
x"00D2",
x"006F",
x"0002",
x"0009",
x"000E",
x"0009",
x"0007",
x"0006",
x"0039",
x"00B5",
x"009A",
x"0034",
x"007E",
x"00BE",
x"00B2",
x"00A2",
x"0084",
x"0063",
x"006F",
x"009A",
x"00B3",
x"00C3",
x"00C5",
x"00CA",
x"00A5",
x"00A1",
x"0057",
x"0052",
x"0014",
x"0004",
x"0001",
x"0005",
x"0007",
x"0008",
x"0006",
x"0002",
x"0004",
x"0007",
x"0008",
x"0008",
x"0007",
x"0003",
x"0005",
x"0003",
x"0002",
x"0005",
x"0014",
x"0022",
x"002F",
x"0051",
x"0054",
x"0058",
x"005C",
x"004A",
x"0038",
x"0036",
x"0044",
x"0061",
x"0080",
x"00AA",
x"00A1",
x"00B1",
x"0078",
x"003D",
x"007C",
x"008F",
x"0079",
x"0047",
x"0045",
x"005E",
x"0063",
x"008F",
x"00B9",
x"00B4",
x"009D",
x"0094",
x"0091",
x"0090",
x"0092",
x"00A0",
x"0098",
x"007B",
x"009A",
x"0094",
x"009A",
x"00A0",
x"0098",
x"008F",
x"0076",
x"007E",
x"0084",
x"0083",
x"0091",
x"0092",
x"0095",
x"0094",
x"0088",
x"008E",
x"008A",
x"0081",
x"0091",
x"009E",
x"008C",
x"0086",
x"0088",
x"0096",
x"0088",
x"007F",
x"007F",
x"0000",
x"0000",
x"0000",
x"0000",
x"00C5",
x"00C5",
x"00C6",
x"00C7",
x"00C5",
x"00C5",
x"00C5",
x"00C4",
x"00C4",
x"00C5",
x"00C4",
x"00C3",
x"00C7",
x"00C8",
x"00C6",
x"00C5",
x"00C5",
x"00C3",
x"00C7",
x"00CC",
x"00BA",
x"0045",
x"0002",
x"0009",
x"0008",
x"0005",
x"0008",
x"005F",
x"00BD",
x"0075",
x"002C",
x"00B7",
x"00CD",
x"00A5",
x"0081",
x"008F",
x"0074",
x"00AA",
x"00C8",
x"00C3",
x"00C1",
x"00C0",
x"00C0",
x"00B3",
x"0081",
x"0072",
x"0098",
x"00A2",
x"0076",
x"003B",
x"0017",
x"0009",
x"0006",
x"000D",
x"0038",
x"0025",
x"000C",
x"0018",
x"0008",
x"000D",
x"0021",
x"0022",
x"002C",
x"0048",
x"0048",
x"0046",
x"0054",
x"003E",
x"0037",
x"0043",
x"004A",
x"005A",
x"006F",
x"0095",
x"00AA",
x"00BF",
x"00D9",
x"00E1",
x"00DD",
x"00AC",
x"00B5",
x"0072",
x"0025",
x"0035",
x"0057",
x"004E",
x"0042",
x"0069",
x"009C",
x"00B7",
x"00B2",
x"00A4",
x"0093",
x"0093",
x"0095",
x"0097",
x"0093",
x"0090",
x"009F",
x"009A",
x"0083",
x"009A",
x"009A",
x"009B",
x"009B",
x"0092",
x"008C",
x"006D",
x"008A",
x"008E",
x"007B",
x"0093",
x"0085",
x"008C",
x"0094",
x"0085",
x"0093",
x"0098",
x"008F",
x"0095",
x"009A",
x"0094",
x"008B",
x"0092",
x"008F",
x"0090",
x"008F",
x"007D",
x"0000",
x"0000",
x"0000",
x"0000",
x"00C4",
x"00C3",
x"00C6",
x"00C7",
x"00C5",
x"00C3",
x"00C5",
x"00C4",
x"00C3",
x"00C5",
x"00C4",
x"00C4",
x"00C6",
x"00C6",
x"00C4",
x"00C3",
x"00C4",
x"00C2",
x"00C5",
x"00C7",
x"00C8",
x"00A9",
x"0040",
x"0004",
x"0009",
x"0008",
x"0008",
x"001A",
x"0064",
x"0087",
x"0067",
x"00C3",
x"00DE",
x"00C5",
x"0056",
x"009A",
x"00B4",
x"00BC",
x"00B9",
x"00B7",
x"00B8",
x"00C7",
x"00C2",
x"00C0",
x"00C6",
x"0092",
x"0082",
x"00C0",
x"00CB",
x"00C1",
x"00A2",
x"002F",
x"0008",
x"0066",
x"009A",
x"005D",
x"005C",
x"0046",
x"0013",
x"0065",
x"007F",
x"0068",
x"0046",
x"002A",
x"001F",
x"0016",
x"0007",
x"0000",
x"0050",
x"009B",
x"00A2",
x"00AA",
x"00AB",
x"00A7",
x"00A4",
x"00AF",
x"00BA",
x"00C1",
x"00C5",
x"009A",
x"00A4",
x"0063",
x"0025",
x"004E",
x"0067",
x"0084",
x"00A1",
x"0096",
x"0091",
x"008C",
x"009D",
x"00A7",
x"0097",
x"0098",
x"0099",
x"0098",
x"0097",
x"0092",
x"00A3",
x"009D",
x"0090",
x"009B",
x"009B",
x"00A0",
x"0094",
x"008F",
x"0095",
x"007E",
x"008B",
x"0083",
x"0078",
x"009A",
x"008F",
x"0089",
x"008C",
x"008A",
x"0099",
x"009F",
x"009D",
x"0093",
x"00A0",
x"0097",
x"0096",
x"009D",
x"008D",
x"0092",
x"0097",
x"0087",
x"0000",
x"0000",
x"0000",
x"0000",
x"00C4",
x"00C3",
x"00C5",
x"00C6",
x"00C4",
x"00C3",
x"00C7",
x"00C3",
x"00C2",
x"00C6",
x"00C3",
x"00C3",
x"00C6",
x"00C6",
x"00C2",
x"00C3",
x"00C3",
x"00C2",
x"00C4",
x"00C6",
x"00C5",
x"00A9",
x"006B",
x"000F",
x"0006",
x"0009",
x"0007",
x"0008",
x"003C",
x"004B",
x"0069",
x"0068",
x"00A6",
x"00BB",
x"005D",
x"0059",
x"0062",
x"0062",
x"0065",
x"0064",
x"0056",
x"0061",
x"009F",
x"00C7",
x"00A5",
x"0040",
x"006B",
x"00C4",
x"00B5",
x"00BB",
x"00C6",
x"0039",
x"0003",
x"001F",
x"0010",
x"0052",
x"00BE",
x"007E",
x"000F",
x"0021",
x"0015",
x"0014",
x"0028",
x"002E",
x"0030",
x"0034",
x"0035",
x"0035",
x"0043",
x"004D",
x"004D",
x"004D",
x"004F",
x"004F",
x"0052",
x"0055",
x"0057",
x"0058",
x"0059",
x"0056",
x"0057",
x"004B",
x"0050",
x"009A",
x"009A",
x"0079",
x"0052",
x"003B",
x"004D",
x"0050",
x"0050",
x"0059",
x"0054",
x"0055",
x"005A",
x"0056",
x"0057",
x"0054",
x"0055",
x"0065",
x"0097",
x"009A",
x"0093",
x"009B",
x"008C",
x"008B",
x"008F",
x"007D",
x"008D",
x"0077",
x"0076",
x"0091",
x"0099",
x"008F",
x"0093",
x"008E",
x"0090",
x"0094",
x"008C",
x"0081",
x"0098",
x"0097",
x"009A",
x"009A",
x"0083",
x"0091",
x"0092",
x"0093",
x"0000",
x"0000",
x"0000",
x"0000",
x"00C5",
x"00C4",
x"00C5",
x"00C6",
x"00C5",
x"00C4",
x"00C6",
x"00C4",
x"00C2",
x"00C4",
x"00C4",
x"00C3",
x"00C8",
x"00C7",
x"00C4",
x"00C4",
x"00C3",
x"00C0",
x"00C3",
x"00C5",
x"00C6",
x"00B6",
x"007A",
x"0030",
x"000D",
x"0008",
x"0004",
x"000B",
x"001C",
x"0037",
x"0060",
x"005E",
x"0042",
x"003A",
x"0038",
x"0038",
x"003D",
x"003F",
x"003D",
x"003F",
x"0044",
x"0048",
x"0035",
x"009B",
x"00A0",
x"0042",
x"006C",
x"00BB",
x"00C7",
x"00C6",
x"00A0",
x"0047",
x"001E",
x"0004",
x"0006",
x"005C",
x"004C",
x"0025",
x"0010",
x"0004",
x"0005",
x"004E",
x"0095",
x"00A2",
x"00A5",
x"00A6",
x"00AC",
x"00B0",
x"00AA",
x"00AA",
x"00AC",
x"00AB",
x"00AE",
x"00AE",
x"00AE",
x"00B1",
x"00B1",
x"00AF",
x"00AF",
x"00B0",
x"00B0",
x"00B0",
x"00B3",
x"009F",
x"0048",
x"004E",
x"0074",
x"0091",
x"00AA",
x"00A7",
x"007F",
x"008B",
x"008C",
x"008B",
x"008F",
x"008C",
x"0087",
x"0086",
x"007A",
x"007B",
x"0094",
x"009B",
x"0098",
x"009E",
x"0097",
x"0093",
x"0083",
x"0074",
x"0093",
x"0072",
x"007C",
x"008C",
x"008C",
x"00A5",
x"0099",
x"0091",
x"0097",
x"0087",
x"0090",
x"008A",
x"008A",
x"008A",
x"008D",
x"0096",
x"008F",
x"008C",
x"008A",
x"008C",
x"0000",
x"0000",
x"0000",
x"0000",
x"00C3",
x"00C3",
x"00C6",
x"00C7",
x"00C5",
x"00C5",
x"00C5",
x"00C3",
x"00C1",
x"00C4",
x"00C3",
x"00C4",
x"00C8",
x"00C8",
x"00C5",
x"00C5",
x"00C1",
x"00C0",
x"00C2",
x"00C4",
x"00C3",
x"00C7",
x"00C4",
x"009F",
x"0063",
x"001D",
x"003A",
x"0050",
x"0024",
x"0043",
x"007E",
x"0064",
x"0043",
x"003C",
x"003F",
x"0071",
x"0057",
x"002D",
x"002F",
x"0036",
x"0032",
x"004F",
x"0030",
x"005D",
x"0085",
x"005A",
x"006D",
x"00D6",
x"00E9",
x"00C0",
x"0092",
x"004B",
x"002B",
x"0009",
x"0011",
x"0054",
x"0061",
x"0061",
x"0026",
x"0007",
x"0011",
x"00B2",
x"00E5",
x"00E6",
x"00E5",
x"00E7",
x"00E8",
x"00EA",
x"00E8",
x"00E7",
x"00E7",
x"00E8",
x"00E6",
x"00E5",
x"00E4",
x"00E5",
x"00E6",
x"00E4",
x"00E3",
x"00E4",
x"00E5",
x"00E6",
x"00E1",
x"00A8",
x"0057",
x"0060",
x"00AA",
x"00D1",
x"00E4",
x"00E3",
x"00CF",
x"00E0",
x"00DE",
x"00E0",
x"00E3",
x"00E2",
x"00E2",
x"00E2",
x"00E1",
x"00C8",
x"009B",
x"009B",
x"009D",
x"009B",
x"0092",
x"0096",
x"0087",
x"0083",
x"009C",
x"0077",
x"007A",
x"0098",
x"0093",
x"009B",
x"009A",
x"0090",
x"0095",
x"009A",
x"0090",
x"0091",
x"0090",
x"0093",
x"008E",
x"0084",
x"0090",
x"008D",
x"0090",
x"008F",
x"0000",
x"0000",
x"0000",
x"0000",
x"00C2",
x"00C3",
x"00C6",
x"00C6",
x"00C5",
x"00C6",
x"00C6",
x"00C3",
x"00C2",
x"00C4",
x"00C4",
x"00C5",
x"00C7",
x"00C8",
x"00C6",
x"00C4",
x"00C1",
x"00C0",
x"00C2",
x"00C5",
x"00C2",
x"00C3",
x"00C6",
x"00C9",
x"00C1",
x"00AD",
x"00B4",
x"0083",
x"0033",
x"004D",
x"006B",
x"0054",
x"005C",
x"004A",
x"005C",
x"007B",
x"003D",
x"0033",
x"0032",
x"0034",
x"0030",
x"0045",
x"002E",
x"0060",
x"007C",
x"00C9",
x"00E4",
x"00F2",
x"00EE",
x"00C9",
x"00A6",
x"003C",
x"0002",
x"000B",
x"0006",
x"005D",
x"00B7",
x"00A7",
x"0018",
x"0004",
x"0008",
x"0049",
x"0070",
x"006C",
x"0061",
x"0076",
x"0083",
x"0094",
x"0094",
x"0092",
x"0091",
x"0093",
x"0094",
x"0095",
x"0094",
x"0095",
x"0099",
x"009B",
x"009C",
x"009A",
x"009F",
x"009B",
x"0097",
x"007E",
x"0069",
x"006B",
x"008F",
x"0098",
x"009C",
x"009B",
x"008D",
x"0099",
x"0094",
x"0096",
x"0096",
x"0092",
x"0091",
x"0091",
x"0094",
x"0093",
x"0097",
x"009E",
x"00A9",
x"009B",
x"0093",
x"0092",
x"0088",
x"0084",
x"0097",
x"007A",
x"0082",
x"008B",
x"008B",
x"009B",
x"009C",
x"0098",
x"008E",
x"0088",
x"0099",
x"0094",
x"008B",
x"0090",
x"008C",
x"0086",
x"008B",
x"0087",
x"009A",
x"0086",
x"0000",
x"0000",
x"0000",
x"0000",
x"00C3",
x"00C3",
x"00C5",
x"00C5",
x"00C5",
x"00C3",
x"00C5",
x"00C4",
x"00C3",
x"00C5",
x"00C3",
x"00C4",
x"00C7",
x"00C7",
x"00C5",
x"00C5",
x"00C4",
x"00C1",
x"00C2",
x"00C4",
x"00C2",
x"00C2",
x"00C4",
x"00C4",
x"00C4",
x"00C8",
x"00C6",
x"007F",
x"003E",
x"0053",
x"0053",
x"0059",
x"00A6",
x"0099",
x"0061",
x"0072",
x"0032",
x"0032",
x"0033",
x"002A",
x"003E",
x"0058",
x"0041",
x"0062",
x"0080",
x"00E5",
x"00EC",
x"00D3",
x"00EC",
x"00E8",
x"00F1",
x"006A",
x"0001",
x"0010",
x"000E",
x"005E",
x"00B8",
x"0087",
x"0049",
x"001D",
x"0009",
x"000C",
x"0009",
x"0007",
x"0048",
x"00AA",
x"00AB",
x"00AB",
x"00A9",
x"00A9",
x"00A9",
x"00A8",
x"00A7",
x"00A8",
x"00A3",
x"009B",
x"00A4",
x"00AD",
x"00BA",
x"00A4",
x"00AE",
x"0078",
x"0068",
x"00B9",
x"00B6",
x"0086",
x"003E",
x"003A",
x"007A",
x"0095",
x"009A",
x"009C",
x"0096",
x"0094",
x"008F",
x"0090",
x"008D",
x"008B",
x"0096",
x"0099",
x"0098",
x"0099",
x"00A5",
x"009A",
x"0096",
x"0096",
x"0085",
x"0089",
x"0096",
x"008E",
x"0091",
x"0085",
x"008A",
x"0095",
x"009A",
x"0091",
x"008F",
x"0087",
x"0097",
x"0090",
x"008A",
x"0091",
x"0088",
x"0084",
x"0085",
x"0088",
x"0080",
x"0078",
x"0000",
x"0000",
x"0000",
x"0000",
x"00C4",
x"00C4",
x"00C5",
x"00C4",
x"00C3",
x"00C3",
x"00C6",
x"00C3",
x"00C0",
x"00C3",
x"00C4",
x"00C4",
x"00C6",
x"00C8",
x"00C6",
x"00C6",
x"00C4",
x"00C2",
x"00C3",
x"00C3",
x"00C3",
x"00C3",
x"00C5",
x"00C3",
x"00C3",
x"00C4",
x"00C4",
x"00B0",
x"0053",
x"0054",
x"0052",
x"006A",
x"00CE",
x"005E",
x"0045",
x"003E",
x"0031",
x"0031",
x"0048",
x"003C",
x"004A",
x"0056",
x"002E",
x"0064",
x"007D",
x"00E2",
x"00F3",
x"00F0",
x"00F4",
x"00EC",
x"00F2",
x"007B",
x"0001",
x"0009",
x"0007",
x"002A",
x"0074",
x"005A",
x"0033",
x"0055",
x"0012",
x"0018",
x"0004",
x"002B",
x"00AB",
x"00B9",
x"00B6",
x"00B3",
x"00B1",
x"00B2",
x"00B2",
x"00B2",
x"00B2",
x"00B1",
x"00A3",
x"009B",
x"00A7",
x"00BC",
x"00C8",
x"00B0",
x"00B2",
x"0084",
x"0066",
x"00CC",
x"00CE",
x"0075",
x"0039",
x"0035",
x"007F",
x"009E",
x"009F",
x"00A0",
x"0099",
x"0095",
x"0091",
x"0092",
x"0094",
x"0090",
x"009D",
x"009A",
x"009E",
x"009B",
x"00A6",
x"00A2",
x"008F",
x"0096",
x"0089",
x"008B",
x"0099",
x"008D",
x"00A4",
x"008F",
x"0087",
x"008C",
x"0093",
x"008B",
x"009C",
x"008C",
x"0093",
x"0082",
x"008B",
x"007C",
x"0082",
x"007F",
x"0087",
x"0096",
x"0085",
x"0090",
x"0000",
x"0000",
x"0000",
x"0000",
x"00C3",
x"00C3",
x"00C4",
x"00C5",
x"00C2",
x"00C2",
x"00C6",
x"00C1",
x"00C1",
x"00C4",
x"00C3",
x"00C4",
x"00C7",
x"00C7",
x"00C5",
x"00C6",
x"00C4",
x"00C2",
x"00C2",
x"00C3",
x"00C2",
x"00C4",
x"00C5",
x"00C2",
x"00C3",
x"00C4",
x"00C4",
x"00BA",
x"0079",
x"005C",
x"0052",
x"006A",
x"00CF",
x"00A1",
x"00B7",
x"0090",
x"004D",
x"0033",
x"0036",
x"0050",
x"006E",
x"0055",
x"0026",
x"0079",
x"0097",
x"00DE",
x"00F6",
x"00FC",
x"00D9",
x"009B",
x"00BB",
x"002F",
x"0008",
x"000B",
x"000A",
x"0007",
x"000A",
x"000B",
x"0010",
x"002A",
x"0010",
x"0008",
x"001E",
x"00A5",
x"00C2",
x"00B6",
x"00B3",
x"00B1",
x"00B0",
x"00B2",
x"00B2",
x"00B2",
x"00B0",
x"00AE",
x"00B1",
x"00AF",
x"00B6",
x"00C9",
x"00D1",
x"00B3",
x"009C",
x"008D",
x"0060",
x"006E",
x"008B",
x"00B1",
x"0055",
x"0054",
x"0086",
x"009C",
x"00A1",
x"009E",
x"0093",
x"008F",
x"0091",
x"008B",
x"0093",
x"0090",
x"0097",
x"0098",
x"009C",
x"009C",
x"00A9",
x"00A6",
x"0096",
x"0095",
x"0088",
x"008D",
x"0094",
x"008D",
x"009D",
x"008C",
x"0087",
x"00A0",
x"0097",
x"008B",
x"0090",
x"0093",
x"00A0",
x"0087",
x"008E",
x"0085",
x"009B",
x"0090",
x"007E",
x"0080",
x"0086",
x"008F",
x"0000",
x"0000",
x"0000",
x"0000",
x"00C3",
x"00C2",
x"00C3",
x"00C4",
x"00C1",
x"00C2",
x"00C4",
x"00C1",
x"00C1",
x"00C3",
x"00C0",
x"00C3",
x"00C7",
x"00C7",
x"00C5",
x"00C5",
x"00C4",
x"00C3",
x"00C2",
x"00C2",
x"00C2",
x"00C3",
x"00C5",
x"00C3",
x"00C1",
x"00C3",
x"00C2",
x"00C3",
x"00B1",
x"0082",
x"0055",
x"005F",
x"00C4",
x"006F",
x"0050",
x"003B",
x"0032",
x"0042",
x"0047",
x"005E",
x"0093",
x"0062",
x"0039",
x"008A",
x"00AA",
x"00E1",
x"00DA",
x"0096",
x"0084",
x"00AB",
x"003B",
x"000F",
x"0012",
x"000A",
x"000C",
x"000B",
x"0006",
x"0007",
x"000E",
x"0020",
x"0032",
x"001B",
x"000A",
x"0045",
x"008B",
x"00B4",
x"00BB",
x"00B5",
x"00B1",
x"00B3",
x"00B3",
x"00AE",
x"0096",
x"006C",
x"0079",
x"0079",
x"007B",
x"00BE",
x"00D4",
x"00BD",
x"0089",
x"00AB",
x"0078",
x"005B",
x"005E",
x"009F",
x"00AD",
x"0072",
x"008A",
x"009B",
x"00A1",
x"009E",
x"0092",
x"008E",
x"0095",
x"008F",
x"0093",
x"008F",
x"0096",
x"009A",
x"009F",
x"0096",
x"00A3",
x"00A2",
x"0093",
x"008E",
x"0095",
x"0099",
x"00A1",
x"009D",
x"0089",
x"008E",
x"008C",
x"0097",
x"009C",
x"0086",
x"0081",
x"008D",
x"0099",
x"008A",
x"0090",
x"0094",
x"009D",
x"0087",
x"0078",
x"0072",
x"0086",
x"0085",
x"0000",
x"0000",
x"0000",
x"0000",
x"00C3",
x"00C3",
x"00C4",
x"00C5",
x"00C1",
x"00C2",
x"00C4",
x"00C2",
x"00C0",
x"00C3",
x"00C1",
x"00C1",
x"00C6",
x"00C6",
x"00C5",
x"00C5",
x"00C4",
x"00C0",
x"00C1",
x"00C2",
x"00C1",
x"00C2",
x"00C3",
x"00C1",
x"00C0",
x"00C1",
x"00C0",
x"00C0",
x"00C5",
x"00C7",
x"0060",
x"0078",
x"00D9",
x"009C",
x"0057",
x"0052",
x"0040",
x"0075",
x"0057",
x"005D",
x"0060",
x"004E",
x"004F",
x"0074",
x"0099",
x"00B5",
x"00C4",
x"00A5",
x"008A",
x"0031",
x"0013",
x"0016",
x"0008",
x"0009",
x"0007",
x"0009",
x"000A",
x"0008",
x"0003",
x"0019",
x"0027",
x"0022",
x"0016",
x"0008",
x"0008",
x"0032",
x"0074",
x"00AB",
x"00BB",
x"00B8",
x"00AA",
x"0074",
x"0066",
x"005C",
x"0072",
x"0076",
x"007B",
x"00BA",
x"00D1",
x"00C8",
x"009C",
x"00AD",
x"0068",
x"004E",
x"0078",
x"007A",
x"008A",
x"00B9",
x"0078",
x"0093",
x"00A1",
x"009D",
x"0093",
x"008F",
x"0094",
x"008B",
x"008D",
x"008E",
x"009A",
x"0096",
x"009A",
x"0095",
x"00A5",
x"009D",
x"008D",
x"0091",
x"0097",
x"009E",
x"009C",
x"008E",
x"0082",
x"0093",
x"0090",
x"0096",
x"0099",
x"0088",
x"008F",
x"0093",
x"0086",
x"0089",
x"008C",
x"0088",
x"0092",
x"008C",
x"0083",
x"0084",
x"0083",
x"0085",
x"0000",
x"0000",
x"0000",
x"0000",
x"00C1",
x"00C1",
x"00C2",
x"00C5",
x"00C1",
x"00C1",
x"00C4",
x"00C1",
x"00BF",
x"00C4",
x"00C1",
x"00C1",
x"00C4",
x"00C4",
x"00C5",
x"00C5",
x"00C3",
x"00C0",
x"00C1",
x"00C1",
x"00C0",
x"00C0",
x"00C2",
x"00C1",
x"00C1",
x"00C1",
x"00C0",
x"00C0",
x"00C2",
x"00C6",
x"0087",
x"0090",
x"0094",
x"0062",
x"006D",
x"0087",
x"0091",
x"009C",
x"0066",
x"003E",
x"0031",
x"0046",
x"002C",
x"0010",
x"0046",
x"0022",
x"0045",
x"002C",
x"0007",
x"0007",
x"0010",
x"0022",
x"002B",
x"0008",
x"0003",
x"0007",
x"000A",
x"0006",
x"002A",
x"0099",
x"007C",
x"0042",
x"0037",
x"002C",
x"001D",
x"000C",
x"0005",
x"0023",
x"006E",
x"00A2",
x"0094",
x"0073",
x"0075",
x"0077",
x"0094",
x"0094",
x"0093",
x"00B8",
x"00B8",
x"00C2",
x"00BB",
x"00AD",
x"0082",
x"0070",
x"0081",
x"007A",
x"0057",
x"00A3",
x"00AF",
x"007D",
x"009B",
x"009E",
x"0092",
x"008E",
x"0092",
x"008A",
x"008C",
x"008D",
x"009C",
x"009A",
x"0096",
x"0099",
x"00A1",
x"0098",
x"0087",
x"008F",
x"009A",
x"009D",
x"00A0",
x"0094",
x"0091",
x"0092",
x"0095",
x"0092",
x"008C",
x"0081",
x"0095",
x"0091",
x"0091",
x"0091",
x"0091",
x"0093",
x"0093",
x"0092",
x"0084",
x"0094",
x"0095",
x"0089",
x"0000",
x"0000",
x"0000",
x"0000",
x"00C0",
x"00C0",
x"00C2",
x"00C3",
x"00C1",
x"00BF",
x"00C5",
x"00C0",
x"00C0",
x"00C4",
x"00C1",
x"00C2",
x"00C4",
x"00C3",
x"00C3",
x"00C5",
x"00C3",
x"00C0",
x"00C0",
x"00C0",
x"00BF",
x"00C0",
x"00C1",
x"00C0",
x"00C0",
x"00C2",
x"00BF",
x"00C0",
x"00C1",
x"00C7",
x"0069",
x"004D",
x"0041",
x"002D",
x"0044",
x"0076",
x"0072",
x"0068",
x"005A",
x"0038",
x"003E",
x"004E",
x"0021",
x"000D",
x"0032",
x"0015",
x"0045",
x"0029",
x"0004",
x"0008",
x"0035",
x"008F",
x"00B6",
x"0074",
x"0030",
x"000D",
x"0004",
x"0037",
x"00A5",
x"00BF",
x"00BF",
x"00BC",
x"00AA",
x"006F",
x"0042",
x"0030",
x"001F",
x"0011",
x"0004",
x"0013",
x"0041",
x"0075",
x"0091",
x"008D",
x"009E",
x"0098",
x"0094",
x"00AF",
x"00AB",
x"00B1",
x"008D",
x"009D",
x"007E",
x"0059",
x"0061",
x"007B",
x"0052",
x"0064",
x"00A1",
x"00BB",
x"0080",
x"0096",
x"0097",
x"008E",
x"0090",
x"008E",
x"0090",
x"0091",
x"0097",
x"0094",
x"009C",
x"0099",
x"00A2",
x"0099",
x"0089",
x"00A0",
x"00A3",
x"0095",
x"009D",
x"009F",
x"0099",
x"0092",
x"0097",
x"0094",
x"008D",
x"007D",
x"008D",
x"0088",
x"008D",
x"008E",
x"0094",
x"0093",
x"009A",
x"0094",
x"007F",
x"009D",
x"0091",
x"008D",
x"0000",
x"0000",
x"0000",
x"0000",
x"00C0",
x"00C0",
x"00C2",
x"00C3",
x"00C0",
x"00C0",
x"00C5",
x"00C1",
x"00C1",
x"00C3",
x"00C1",
x"00C1",
x"00C3",
x"00C4",
x"00C3",
x"00C4",
x"00C2",
x"00BF",
x"00C0",
x"00C1",
x"00C0",
x"00C0",
x"00C2",
x"00C0",
x"00BF",
x"00C0",
x"00BF",
x"00BF",
x"00C1",
x"00C6",
x"007D",
x"0046",
x"0088",
x"0093",
x"0091",
x"009C",
x"009D",
x"00B3",
x"009E",
x"0087",
x"005D",
x"0038",
x"001A",
x"0007",
x"002B",
x"0018",
x"0039",
x"002C",
x"0010",
x"004D",
x"00B2",
x"00BE",
x"00BA",
x"00C1",
x"00BA",
x"0088",
x"006E",
x"00A8",
x"00BA",
x"00B5",
x"00B6",
x"00B7",
x"00BA",
x"00C0",
x"00B6",
x"007F",
x"004B",
x"0039",
x"0029",
x"0018",
x"0008",
x"000A",
x"0033",
x"0069",
x"0099",
x"00A6",
x"009A",
x"0089",
x"009B",
x"00AE",
x"00A3",
x"00A9",
x"0086",
x"005C",
x"0059",
x"0074",
x"0065",
x"0065",
x"0083",
x"00AA",
x"00BB",
x"0080",
x"0084",
x"008B",
x"008F",
x"0090",
x"0090",
x"008F",
x"0098",
x"0099",
x"009A",
x"0095",
x"009B",
x"009F",
x"0097",
x"009D",
x"009D",
x"0091",
x"009D",
x"009F",
x"0098",
x"0097",
x"008D",
x"0096",
x"0094",
x"0081",
x"008D",
x"0090",
x"008C",
x"0094",
x"0092",
x"0090",
x"009B",
x"00A0",
x"008D",
x"0095",
x"009D",
x"0099",
x"0000",
x"0000",
x"0000",
x"0000",
x"00BF",
x"00BF",
x"00C2",
x"00C3",
x"00C0",
x"00C2",
x"00C5",
x"00C1",
x"00C1",
x"00C2",
x"00C0",
x"00BF",
x"00C3",
x"00C4",
x"00C2",
x"00C2",
x"00C3",
x"00C0",
x"00C0",
x"00C0",
x"00C0",
x"00C2",
x"00C3",
x"00C0",
x"00BF",
x"00BF",
x"00BF",
x"00BE",
x"00C0",
x"00C0",
x"00C3",
x"00AA",
x"00B9",
x"0081",
x"0057",
x"008C",
x"0084",
x"00B2",
x"0077",
x"0073",
x"0072",
x"005F",
x"002E",
x"0000",
x"0035",
x"004B",
x"0067",
x"0081",
x"0089",
x"00B9",
x"00BA",
x"00B7",
x"00B6",
x"00B7",
x"00B9",
x"00BB",
x"00BE",
x"00B8",
x"00B4",
x"00B5",
x"00B5",
x"00B5",
x"00B6",
x"00B7",
x"00B8",
x"00BC",
x"00B9",
x"0097",
x"005E",
x"003A",
x"0029",
x"001C",
x"000A",
x"0003",
x"0022",
x"0063",
x"009C",
x"00AC",
x"00A6",
x"00AD",
x"008C",
x"00A7",
x"007E",
x"0057",
x"004F",
x"0076",
x"0094",
x"0079",
x"008D",
x"0099",
x"00A9",
x"00BF",
x"0078",
x"007D",
x"008D",
x"008C",
x"0090",
x"008B",
x"009A",
x"009E",
x"009B",
x"0092",
x"009B",
x"0099",
x"0094",
x"009C",
x"0091",
x"008E",
x"009A",
x"0098",
x"0099",
x"009F",
x"0098",
x"009A",
x"008B",
x"0084",
x"0095",
x"008E",
x"0085",
x"008C",
x"0099",
x"0098",
x"0096",
x"0091",
x"0089",
x"0092",
x"008F",
x"0083",
x"0000",
x"0000",
x"0000",
x"0000",
x"00C0",
x"00C0",
x"00C2",
x"00C2",
x"00C2",
x"00C3",
x"00C4",
x"00C1",
x"00BF",
x"00C2",
x"00BF",
x"00BF",
x"00C1",
x"00C1",
x"00C3",
x"00C2",
x"00C1",
x"00C0",
x"00C0",
x"00C1",
x"00BF",
x"00C1",
x"00C2",
x"00C0",
x"00BF",
x"00BF",
x"00BE",
x"00BE",
x"00C0",
x"00BF",
x"00BE",
x"00B0",
x"00CE",
x"0086",
x"005A",
x"007C",
x"0073",
x"00D7",
x"005E",
x"006E",
x"00CC",
x"00C3",
x"008E",
x"005F",
x"009A",
x"00B5",
x"00BD",
x"00C1",
x"00BE",
x"00B8",
x"00B7",
x"00B6",
x"00B5",
x"00B5",
x"00B5",
x"00B5",
x"00B6",
x"00B5",
x"00B5",
x"00B4",
x"00B5",
x"00B5",
x"00B4",
x"00B7",
x"00B6",
x"00B6",
x"00B7",
x"00B9",
x"00C0",
x"00AE",
x"0072",
x"0041",
x"0026",
x"001E",
x"0013",
x"0004",
x"0019",
x"0055",
x"0075",
x"009E",
x"008F",
x"00A3",
x"0087",
x"006A",
x"0063",
x"006F",
x"0089",
x"0087",
x"0098",
x"009C",
x"009A",
x"00AA",
x"00BB",
x"007D",
x"007F",
x"008E",
x"0087",
x"0087",
x"0098",
x"009A",
x"0093",
x"0090",
x"0094",
x"0099",
x"0091",
x"009C",
x"0092",
x"0099",
x"009F",
x"009F",
x"009C",
x"0098",
x"00A0",
x"00A4",
x"0089",
x"0092",
x"0093",
x"0086",
x"008D",
x"008E",
x"0092",
x"009A",
x"009F",
x"0098",
x"0078",
x"0085",
x"0094",
x"008F",
x"0000",
x"0000",
x"0000",
x"0000",
x"00C0",
x"00C0",
x"00C1",
x"00C1",
x"00C0",
x"00C2",
x"00C3",
x"00C0",
x"00C0",
x"00C1",
x"00BF",
x"00BF",
x"00C0",
x"00C0",
x"00C1",
x"00C3",
x"00C1",
x"00C0",
x"00C0",
x"00C0",
x"00BF",
x"00BF",
x"00C1",
x"00C0",
x"00BE",
x"00BF",
x"00BD",
x"00BF",
x"00C0",
x"00BF",
x"00BD",
x"00B6",
x"00D7",
x"008F",
x"0072",
x"00A3",
x"00AE",
x"00DC",
x"0080",
x"0076",
x"00BF",
x"00BA",
x"00BD",
x"00C0",
x"00BC",
x"00B7",
x"00B7",
x"00B7",
x"00B6",
x"00B6",
x"00B5",
x"00B6",
x"00B4",
x"00B5",
x"00B3",
x"00B4",
x"00B4",
x"00B5",
x"00B3",
x"00B2",
x"00B4",
x"00B3",
x"00B4",
x"00B5",
x"00B4",
x"00B5",
x"00B4",
x"00B3",
x"00C1",
x"00D0",
x"00CB",
x"00B1",
x"007D",
x"0049",
x"0032",
x"0026",
x"0018",
x"0006",
x"0009",
x"0030",
x"0069",
x"0093",
x"009E",
x"0091",
x"007D",
x"0053",
x"0064",
x"007C",
x"008E",
x"009C",
x"00A2",
x"009C",
x"009A",
x"00B9",
x"0082",
x"0081",
x"0087",
x"008C",
x"009D",
x"0096",
x"0097",
x"0098",
x"0092",
x"009B",
x"008E",
x"0096",
x"008D",
x"009C",
x"00A0",
x"009C",
x"00A0",
x"0093",
x"009D",
x"00A1",
x"008F",
x"0086",
x"008A",
x"0080",
x"0096",
x"009F",
x"008C",
x"008F",
x"0091",
x"008D",
x"007E",
x"0087",
x"009A",
x"0090",
x"0000",
x"0000",
x"0000",
x"0000",
x"00BF",
x"00BF",
x"00C0",
x"00C1",
x"00C0",
x"00C1",
x"00C2",
x"00BF",
x"00BF",
x"00BF",
x"00BD",
x"00BF",
x"00BF",
x"00C0",
x"00BF",
x"00C1",
x"00C1",
x"00C0",
x"00BF",
x"00BF",
x"00BF",
x"00BF",
x"00C1",
x"00BF",
x"00BE",
x"00C0",
x"00BE",
x"00BE",
x"00BE",
x"00BE",
x"00BE",
x"00AF",
x"00CE",
x"008A",
x"0098",
x"00C4",
x"00B6",
x"00D7",
x"0072",
x"0070",
x"00BF",
x"00BA",
x"00B8",
x"00B7",
x"00B7",
x"00B6",
x"00B5",
x"00B6",
x"00B6",
x"00B5",
x"00B5",
x"00B6",
x"00B2",
x"00B4",
x"00B4",
x"00B4",
x"00B3",
x"00B3",
x"00B2",
x"00B2",
x"00B4",
x"00B3",
x"00B4",
x"00B4",
x"00B4",
x"00B4",
x"00B1",
x"00B5",
x"00C8",
x"00C9",
x"00C6",
x"00C2",
x"00BE",
x"00B4",
x"00A0",
x"0069",
x"003E",
x"0027",
x"0021",
x"000B",
x"0002",
x"001E",
x"0057",
x"0089",
x"0091",
x"007D",
x"0082",
x"0076",
x"008F",
x"009D",
x"009F",
x"009D",
x"0087",
x"0090",
x"00BB",
x"0089",
x"0076",
x"008A",
x"009D",
x"009C",
x"009B",
x"0090",
x"0095",
x"009E",
x"0092",
x"0097",
x"009B",
x"009A",
x"0097",
x"009D",
x"009E",
x"0090",
x"008E",
x"00A4",
x"0089",
x"0086",
x"008F",
x"0080",
x"008E",
x"0092",
x"0098",
x"008F",
x"008D",
x"0092",
x"0089",
x"0085",
x"0096",
x"0097",
x"0000",
x"0000",
x"0000",
x"0000",
x"00BE",
x"00BE",
x"00C0",
x"00BF",
x"00BF",
x"00C0",
x"00C0",
x"00BD",
x"00BF",
x"00BF",
x"00BD",
x"00BF",
x"00BF",
x"00BE",
x"00BF",
x"00C1",
x"00BF",
x"00BE",
x"00BE",
x"00BE",
x"00BD",
x"00BF",
x"00C0",
x"00BE",
x"00BE",
x"00BF",
x"00BE",
x"00BD",
x"00BE",
x"00BE",
x"00BD",
x"00BD",
x"00BD",
x"00B8",
x"00BD",
x"00BF",
x"00B0",
x"00D8",
x"0071",
x"006A",
x"00BF",
x"00BA",
x"00B6",
x"00B7",
x"00B7",
x"00B5",
x"00B4",
x"00B4",
x"00B4",
x"00B2",
x"00B2",
x"00B3",
x"00B2",
x"00B3",
x"00B4",
x"00B3",
x"00B2",
x"00B2",
x"00B2",
x"00B2",
x"00B2",
x"00B3",
x"00B3",
x"00B3",
x"00B2",
x"00B2",
x"00B2",
x"00B5",
x"00CB",
x"00CD",
x"00C9",
x"00C5",
x"00B9",
x"00BD",
x"00C8",
x"00C1",
x"00AE",
x"0079",
x"0037",
x"0022",
x"001C",
x"000D",
x"0004",
x"001B",
x"0042",
x"006C",
x"008A",
x"0085",
x"0095",
x"009D",
x"009C",
x"0099",
x"008C",
x"0088",
x"0092",
x"00BC",
x"0081",
x"0073",
x"00A1",
x"00A0",
x"009A",
x"0095",
x"0092",
x"0098",
x"0090",
x"0097",
x"0098",
x"0091",
x"0094",
x"0097",
x"00A1",
x"00A2",
x"009C",
x"0099",
x"0088",
x"008C",
x"008F",
x"008C",
x"0096",
x"008D",
x"0092",
x"008C",
x"0096",
x"0094",
x"009D",
x"007A",
x"0075",
x"0090",
x"0000",
x"0000",
x"0000",
x"0000",
x"00BD",
x"00BE",
x"00C0",
x"00BF",
x"00BD",
x"00BF",
x"00C1",
x"00BD",
x"00BC",
x"00BE",
x"00BC",
x"00BC",
x"00BF",
x"00BE",
x"00BE",
x"00C0",
x"00BF",
x"00BD",
x"00BF",
x"00BD",
x"00BB",
x"00BD",
x"00BF",
x"00BE",
x"00BE",
x"00BF",
x"00BC",
x"00BD",
x"00BD",
x"00BE",
x"00BD",
x"00BF",
x"00BC",
x"00BC",
x"00BC",
x"00BB",
x"008B",
x"0070",
x"0030",
x"005C",
x"00BE",
x"00B8",
x"00B5",
x"00B5",
x"00B5",
x"00B4",
x"00B5",
x"00B5",
x"00B4",
x"00B1",
x"00B2",
x"00B3",
x"00B2",
x"00B4",
x"00B2",
x"00B2",
x"00B2",
x"00B2",
x"00B1",
x"00B2",
x"00B2",
x"00B1",
x"00B2",
x"00B2",
x"00B2",
x"00B2",
x"00B1",
x"00B2",
x"00CA",
x"00D3",
x"00CB",
x"00C7",
x"00BB",
x"00BC",
x"009D",
x"00AC",
x"00C5",
x"00C7",
x"009D",
x"0081",
x"0042",
x"0029",
x"0022",
x"0015",
x"0004",
x"000A",
x"0031",
x"0062",
x"0095",
x"00A5",
x"00A6",
x"0099",
x"008D",
x"0088",
x"0085",
x"008F",
x"00BB",
x"0090",
x"0084",
x"009F",
x"0099",
x"0099",
x"008A",
x"009B",
x"0096",
x"0097",
x"0094",
x"0097",
x"009C",
x"0097",
x"00A3",
x"009D",
x"0090",
x"009B",
x"0095",
x"0093",
x"00A3",
x"0094",
x"0095",
x"0090",
x"009A",
x"008B",
x"008C",
x"0090",
x"009D",
x"008C",
x"007E",
x"0086",
x"0000",
x"0000",
x"0000",
x"0000",
x"00BE",
x"00BE",
x"00BE",
x"00BE",
x"00BE",
x"00BF",
x"00C0",
x"00BD",
x"00BD",
x"00BF",
x"00BC",
x"00BD",
x"00BE",
x"00BE",
x"00BF",
x"00BF",
x"00BE",
x"00BD",
x"00BE",
x"00BC",
x"00BC",
x"00BC",
x"00BE",
x"00BD",
x"00BD",
x"00BE",
x"00BC",
x"00BB",
x"00BC",
x"00BD",
x"00BC",
x"00BD",
x"00BC",
x"00BB",
x"00BB",
x"00C2",
x"0080",
x"003D",
x"0009",
x"0052",
x"00C0",
x"00B8",
x"00B5",
x"00B6",
x"00B5",
x"00B4",
x"00B5",
x"00B5",
x"00B4",
x"00B2",
x"00B2",
x"00B2",
x"00B2",
x"00B3",
x"00B2",
x"00B2",
x"00B2",
x"00B1",
x"00B1",
x"00B1",
x"00B1",
x"00B1",
x"00B2",
x"00B2",
x"00B2",
x"00B1",
x"00B2",
x"00B0",
x"00C2",
x"00D5",
x"00CC",
x"00C7",
x"00BF",
x"00B5",
x"00A3",
x"00B7",
x"00C2",
x"00BC",
x"00AF",
x"00B5",
x"0075",
x"0068",
x"0042",
x"0024",
x"0024",
x"0018",
x"0005",
x"0008",
x"0027",
x"005B",
x"009B",
x"009E",
x"0090",
x"0089",
x"0087",
x"008A",
x"008B",
x"00AE",
x"0096",
x"007E",
x"0097",
x"0097",
x"0096",
x"00A2",
x"0094",
x"0097",
x"0094",
x"008D",
x"0093",
x"0091",
x"00A0",
x"0089",
x"0093",
x"009A",
x"0091",
x"0083",
x"0090",
x"0083",
x"0098",
x"0095",
x"009D",
x"0093",
x"0092",
x"0091",
x"0091",
x"008D",
x"008C",
x"00A0",
x"0000",
x"0000",
x"0000",
x"0000",
x"00BD",
x"00BD",
x"00BF",
x"00BE",
x"00BD",
x"00BF",
x"00BE",
x"00BB",
x"00BC",
x"00BC",
x"00BB",
x"00BE",
x"00BF",
x"00BE",
x"00BF",
x"00BF",
x"00BE",
x"00BC",
x"00BE",
x"00BB",
x"00BA",
x"00BD",
x"00BF",
x"00BD",
x"00BE",
x"00BD",
x"00BA",
x"00BB",
x"00BC",
x"00BB",
x"00BC",
x"00BC",
x"00BC",
x"00BA",
x"00BA",
x"00BD",
x"00A7",
x"009A",
x"0076",
x"0091",
x"00BB",
x"00B6",
x"00B4",
x"00B6",
x"00B6",
x"00B4",
x"00B4",
x"00B5",
x"00B4",
x"00B2",
x"00B2",
x"00B1",
x"00B1",
x"00B2",
x"00B2",
x"00B1",
x"00B2",
x"00B2",
x"00B0",
x"00B1",
x"00B1",
x"00B2",
x"00B1",
x"00B2",
x"00B2",
x"00B2",
x"00B1",
x"00B0",
x"00B6",
x"00D0",
x"00D0",
x"00C8",
x"00C4",
x"00BC",
x"00B4",
x"00BB",
x"00C3",
x"00BC",
x"00AE",
x"00A2",
x"0038",
x"0037",
x"003A",
x"002E",
x"002F",
x"002A",
x"001F",
x"001C",
x"000B",
x"0004",
x"001C",
x"0046",
x"0073",
x"008E",
x"008B",
x"0088",
x"0083",
x"0086",
x"00B9",
x"0095",
x"007A",
x"0098",
x"0099",
x"0097",
x"0090",
x"008E",
x"0090",
x"0084",
x"0099",
x"00A2",
x"00A1",
x"0091",
x"0092",
x"0097",
x"0095",
x"0092",
x"0097",
x"0089",
x"0083",
x"008F",
x"00A2",
x"008F",
x"0088",
x"0090",
x"009F",
x"0094",
x"0086",
x"0091",
x"0000",
x"0000",
x"0000",
x"0000",
x"00BC",
x"00BD",
x"00BE",
x"00BE",
x"00BC",
x"00BE",
x"00BF",
x"00BB",
x"00BB",
x"00BD",
x"00BA",
x"00BC",
x"00BE",
x"00BD",
x"00BE",
x"00BF",
x"00BD",
x"00BD",
x"00BE",
x"00BD",
x"00BA",
x"00BC",
x"00BE",
x"00BD",
x"00BE",
x"00BD",
x"00BA",
x"00BA",
x"00BB",
x"00BB",
x"00BC",
x"00BC",
x"00BA",
x"00BA",
x"00BA",
x"00B8",
x"00BC",
x"00C0",
x"00C2",
x"00BE",
x"00B8",
x"00B8",
x"00B6",
x"00B5",
x"00B6",
x"00B4",
x"00B3",
x"00B5",
x"00B5",
x"00B2",
x"00B2",
x"00B1",
x"00B1",
x"00B3",
x"00B3",
x"00B2",
x"00B2",
x"00B2",
x"00B1",
x"00B0",
x"00B1",
x"00B2",
x"00B3",
x"00B3",
x"00B3",
x"00B3",
x"00B1",
x"00B1",
x"00AF",
x"00BD",
x"00CD",
x"00CA",
x"00C5",
x"00C4",
x"00BF",
x"00C0",
x"00C2",
x"00B9",
x"00A9",
x"00B6",
x"008F",
x"0098",
x"0098",
x"0098",
x"0095",
x"0091",
x"005C",
x"0038",
x"0024",
x"001C",
x"000F",
x"0003",
x"000E",
x"0034",
x"0064",
x"008A",
x"0091",
x"0088",
x"009C",
x"00BA",
x"0095",
x"0078",
x"0092",
x"0092",
x"0097",
x"009A",
x"0093",
x"0081",
x"0097",
x"00A1",
x"009D",
x"0093",
x"009A",
x"00A2",
x"009C",
x"0091",
x"0094",
x"0099",
x"007F",
x"0087",
x"009B",
x"0093",
x"0085",
x"0093",
x"0096",
x"008B",
x"008F",
x"0084",
x"0000",
x"0000",
x"0000",
x"0000",
x"00BB",
x"00BC",
x"00BD",
x"00BD",
x"00BB",
x"00BD",
x"00BD",
x"00BA",
x"00BB",
x"00BC",
x"00BA",
x"00BB",
x"00BC",
x"00BB",
x"00BD",
x"00BF",
x"00BD",
x"00BD",
x"00BD",
x"00BC",
x"00BA",
x"00BB",
x"00BE",
x"00BD",
x"00BC",
x"00BD",
x"00BC",
x"00BC",
x"00BC",
x"00BA",
x"00BB",
x"00BB",
x"00BA",
x"00BB",
x"00BA",
x"00B9",
x"00B8",
x"00BA",
x"00BB",
x"00B9",
x"00B7",
x"00B8",
x"00B5",
x"00B6",
x"00B7",
x"00B5",
x"00B5",
x"00B6",
x"00B6",
x"00B3",
x"00B3",
x"00B2",
x"00B1",
x"00B2",
x"00B3",
x"00B1",
x"00B2",
x"00B2",
x"00B1",
x"00B2",
x"00B2",
x"00B3",
x"00B3",
x"00B2",
x"00B2",
x"00B1",
x"00B2",
x"00B1",
x"00AF",
x"00B0",
x"00BE",
x"00C9",
x"00C8",
x"00C9",
x"00C7",
x"00C0",
x"00C1",
x"00BB",
x"00AB",
x"009B",
x"0038",
x"0042",
x"0059",
x"0062",
x"0057",
x"0051",
x"0064",
x"0085",
x"0079",
x"004E",
x"002C",
x"001E",
x"0013",
x"0006",
x"0009",
x"0025",
x"0054",
x"007C",
x"009E",
x"009E",
x"00B8",
x"0098",
x"0075",
x"0092",
x"0092",
x"0096",
x"008B",
x"008E",
x"0092",
x"0091",
x"00A1",
x"0096",
x"0097",
x"0099",
x"0098",
x"0087",
x"0092",
x"008C",
x"007A",
x"0087",
x"0097",
x"0099",
x"008B",
x"009F",
x"009F",
x"0092",
x"007D",
x"0087",
x"0000",
x"0000",
x"0000",
x"0000",
x"00BC",
x"00BC",
x"00BD",
x"00BB",
x"00BB",
x"00BC",
x"00BE",
x"00BA",
x"00BA",
x"00BA",
x"00B9",
x"00BC",
x"00BC",
x"00BA",
x"00BD",
x"00BF",
x"00BF",
x"00BC",
x"00BC",
x"00BA",
x"00B9",
x"00BA",
x"00BD",
x"00BD",
x"00BC",
x"00BB",
x"00BA",
x"00BC",
x"00BB",
x"00BA",
x"00BB",
x"00BC",
x"00BA",
x"00B9",
x"00B8",
x"00B8",
x"00B8",
x"00BA",
x"00BA",
x"00B7",
x"00B8",
x"00B7",
x"00B5",
x"00B6",
x"00B5",
x"00B5",
x"00B5",
x"00B6",
x"00B4",
x"00B3",
x"00B3",
x"00B2",
x"00B1",
x"00B2",
x"00B1",
x"00AF",
x"00B0",
x"00B1",
x"00B1",
x"00B1",
x"00B2",
x"00B1",
x"00B2",
x"00B1",
x"00B1",
x"00B1",
x"00B1",
x"00B1",
x"00AF",
x"00AF",
x"00AE",
x"00BF",
x"00CE",
x"00CD",
x"00C9",
x"00BB",
x"00C3",
x"00BD",
x"00A5",
x"00AE",
x"006C",
x"0068",
x"0070",
x"006C",
x"005B",
x"005C",
x"007A",
x"0082",
x"009C",
x"00A5",
x"0091",
x"005A",
x"0030",
x"0021",
x"0019",
x"000A",
x"0006",
x"0014",
x"0047",
x"007F",
x"0096",
x"00B4",
x"0098",
x"0079",
x"0090",
x"008C",
x"008C",
x"0093",
x"0099",
x"009D",
x"0096",
x"0093",
x"009A",
x"0093",
x"008D",
x"0087",
x"008F",
x"008F",
x"007F",
x"008E",
x"008B",
x"0092",
x"0097",
x"0098",
x"008F",
x"009B",
x"0092",
x"0090",
x"0000",
x"0000",
x"0000",
x"0000",
x"00BC",
x"00BC",
x"00BC",
x"00BB",
x"00BA",
x"00BD",
x"00BD",
x"00BA",
x"00BA",
x"00BB",
x"00B9",
x"00B9",
x"00BC",
x"00B9",
x"00BD",
x"00BF",
x"00BD",
x"00BA",
x"00BA",
x"00BA",
x"00BB",
x"00BB",
x"00BC",
x"00BB",
x"00BD",
x"00BC",
x"00B9",
x"00B9",
x"00BA",
x"00BB",
x"00B9",
x"00BB",
x"00B9",
x"00B9",
x"00BA",
x"00B8",
x"00B9",
x"00BB",
x"00BA",
x"00B7",
x"00B8",
x"00B7",
x"00B5",
x"00B6",
x"00B6",
x"00B4",
x"00B6",
x"00B7",
x"00B4",
x"00B3",
x"00B3",
x"00B1",
x"00B1",
x"00B1",
x"00B1",
x"00B1",
x"00B1",
x"00B0",
x"00B0",
x"00B1",
x"00B2",
x"00B0",
x"00B1",
x"00B1",
x"00B0",
x"00B1",
x"00B2",
x"00B0",
x"00AF",
x"00B1",
x"00BB",
x"00A8",
x"00C5",
x"00D3",
x"00C9",
x"00BA",
x"00BE",
x"00BA",
x"00A8",
x"009F",
x"0053",
x"005D",
x"0067",
x"0069",
x"0060",
x"006A",
x"008E",
x"007B",
x"0095",
x"009F",
x"00A2",
x"00A1",
x"0088",
x"0068",
x"0039",
x"0022",
x"0019",
x"000E",
x"0005",
x"0010",
x"003A",
x"0064",
x"00B0",
x"00D4",
x"00A8",
x"0093",
x"0092",
x"008A",
x"009F",
x"00A1",
x"009C",
x"0090",
x"0091",
x"0092",
x"0095",
x"0099",
x"009B",
x"008A",
x"0086",
x"0090",
x"0090",
x"008B",
x"0093",
x"009B",
x"0095",
x"008F",
x"0090",
x"008A",
x"0000",
x"0000",
x"0000",
x"0000",
x"00BA",
x"00B9",
x"00BA",
x"00B9",
x"00B9",
x"00BC",
x"00BC",
x"00BA",
x"00B9",
x"00B9",
x"00B8",
x"00B9",
x"00BA",
x"00B8",
x"00BC",
x"00BD",
x"00BC",
x"00BA",
x"00B9",
x"00BA",
x"00B9",
x"00BC",
x"00BC",
x"00BB",
x"00BB",
x"00BA",
x"00B9",
x"00BA",
x"00BA",
x"00B9",
x"00B9",
x"00BB",
x"00B9",
x"00B9",
x"00BA",
x"00B8",
x"00B7",
x"00B9",
x"00B8",
x"00B7",
x"00B7",
x"00B7",
x"00B5",
x"00B6",
x"00B7",
x"00B5",
x"00B5",
x"00B6",
x"00B4",
x"00B4",
x"00B4",
x"00B1",
x"00B1",
x"00B2",
x"00B2",
x"00B1",
x"00AF",
x"00B0",
x"00AF",
x"00B1",
x"00B1",
x"00B1",
x"00B1",
x"00B1",
x"00B0",
x"00B1",
x"00B1",
x"00B1",
x"00B0",
x"00B0",
x"00BB",
x"00A3",
x"00BB",
x"00D3",
x"00CC",
x"00BC",
x"00B8",
x"00B7",
x"00A8",
x"009B",
x"0042",
x"0040",
x"004F",
x"005A",
x"0054",
x"005B",
x"0087",
x"0072",
x"0093",
x"009C",
x"009C",
x"0099",
x"008E",
x"0093",
x"0085",
x"006D",
x"0042",
x"002B",
x"0018",
x"000E",
x"0008",
x"0006",
x"0054",
x"00B1",
x"0093",
x"008B",
x"008B",
x"008C",
x"009D",
x"00A5",
x"00A3",
x"009A",
x"0097",
x"008D",
x"0090",
x"0094",
x"00A4",
x"008A",
x"0079",
x"0086",
x"0094",
x"008E",
x"0090",
x"00A1",
x"009A",
x"0085",
x"0088",
x"009A",
x"0000",
x"0000",
x"0000",
x"0000",
x"00B8",
x"00B8",
x"00B9",
x"00B9",
x"00B8",
x"00BA",
x"00BB",
x"00BB",
x"00BA",
x"00B9",
x"00B7",
x"00B8",
x"00B8",
x"00B7",
x"00BA",
x"00BC",
x"00BA",
x"00B8",
x"00B9",
x"00B9",
x"00B8",
x"00B9",
x"00BA",
x"00BA",
x"00BA",
x"00BC",
x"00B8",
x"00B7",
x"00B8",
x"00B8",
x"00B7",
x"00BA",
x"00B9",
x"00B8",
x"00B8",
x"00B8",
x"00B7",
x"00B8",
x"00B9",
x"00B8",
x"00B7",
x"00B7",
x"00B4",
x"00B5",
x"00B7",
x"00B6",
x"00B4",
x"00B6",
x"00B4",
x"00B4",
x"00B4",
x"00B2",
x"00B1",
x"00B1",
x"00B2",
x"00B1",
x"00B0",
x"00AF",
x"00AE",
x"00B0",
x"00B1",
x"00B1",
x"00B0",
x"00B1",
x"00B0",
x"00AF",
x"00B0",
x"00B0",
x"00AF",
x"00B0",
x"00B9",
x"00A3",
x"00B2",
x"00CB",
x"00CE",
x"00C1",
x"00BC",
x"00B6",
x"00A5",
x"00A9",
x"0099",
x"00B2",
x"00A6",
x"0090",
x"0079",
x"008F",
x"0099",
x"006C",
x"008F",
x"009D",
x"009E",
x"0097",
x"008A",
x"008A",
x"0083",
x"008C",
x"008F",
x"0082",
x"0055",
x"002F",
x"001C",
x"001D",
x"008F",
x"005E",
x"0015",
x"0048",
x"0073",
x"00A1",
x"00A6",
x"009E",
x"0092",
x"0092",
x"0096",
x"0090",
x"009A",
x"0093",
x"00A4",
x"0093",
x"007C",
x"0084",
x"008B",
x"0085",
x"008B",
x"009E",
x"0093",
x"008F",
x"008A",
x"0092",
x"0000",
x"0000",
x"0000",
x"0000",
x"00B8",
x"00B8",
x"00B8",
x"00B9",
x"00B7",
x"00B8",
x"00B8",
x"00B7",
x"00B9",
x"00B8",
x"00B6",
x"00B6",
x"00B8",
x"00B7",
x"00B8",
x"00BA",
x"00B9",
x"00BB",
x"00BB",
x"00B8",
x"00B8",
x"00B8",
x"00B8",
x"00B8",
x"00B9",
x"00B9",
x"00B8",
x"00B6",
x"00B8",
x"00B8",
x"00B6",
x"00B9",
x"00B8",
x"00B6",
x"00B8",
x"00B7",
x"00B7",
x"00B8",
x"00B7",
x"00B6",
x"00B6",
x"00B6",
x"00B4",
x"00B5",
x"00B5",
x"00B5",
x"00B4",
x"00B4",
x"00B3",
x"00B2",
x"00B1",
x"00B1",
x"00B0",
x"00B0",
x"00B1",
x"00B0",
x"00B0",
x"00B0",
x"00AE",
x"00AF",
x"00AF",
x"00AF",
x"00B0",
x"00B0",
x"00AF",
x"00AE",
x"00B0",
x"00B0",
x"00AF",
x"00AE",
x"00B7",
x"00A1",
x"00AA",
x"00AE",
x"00C6",
x"00BF",
x"00B8",
x"00B5",
x"00A5",
x"008C",
x"0053",
x"0074",
x"0067",
x"0065",
x"006B",
x"0074",
x"0083",
x"0071",
x"0092",
x"009B",
x"009A",
x"0093",
x"008B",
x"008C",
x"007E",
x"0086",
x"0089",
x"0092",
x"00A2",
x"0096",
x"0060",
x"006D",
x"00E6",
x"006B",
x"0006",
x"0005",
x"000E",
x"0047",
x"007C",
x"0090",
x"0098",
x"009C",
x"008E",
x"0085",
x"008E",
x"0091",
x"0095",
x"008F",
x"0086",
x"008D",
x"008A",
x"0089",
x"008A",
x"0085",
x"0093",
x"008E",
x"0086",
x"0081",
x"0000",
x"0000",
x"0000",
x"0000",
x"00B7",
x"00B7",
x"00B7",
x"00B7",
x"00B8",
x"00B7",
x"00B8",
x"00B5",
x"00B6",
x"00B8",
x"00B5",
x"00B7",
x"00B9",
x"00B7",
x"00B9",
x"00BA",
x"00B8",
x"00BA",
x"00B9",
x"00B8",
x"00B7",
x"00B9",
x"00B9",
x"00B8",
x"00B9",
x"00B8",
x"00B8",
x"00B7",
x"00B8",
x"00B7",
x"00B7",
x"00B9",
x"00B7",
x"00B7",
x"00B8",
x"00B7",
x"00B6",
x"00B7",
x"00B7",
x"00B6",
x"00B6",
x"00B5",
x"00B4",
x"00B4",
x"00B4",
x"00B5",
x"00B3",
x"00B4",
x"00B3",
x"00B2",
x"00B2",
x"00B1",
x"00B0",
x"00B1",
x"00B1",
x"00B0",
x"00B0",
x"00B0",
x"00AE",
x"00AF",
x"00B0",
x"00B0",
x"00AF",
x"00B0",
x"00AF",
x"00AF",
x"00AE",
x"00AF",
x"00AD",
x"00B0",
x"00B8",
x"009F",
x"00AB",
x"00A0",
x"00A5",
x"00C0",
x"00BF",
x"00AF",
x"009A",
x"00B5",
x"00AD",
x"00AC",
x"0082",
x"0049",
x"0043",
x"0049",
x"0059",
x"0074",
x"0093",
x"009E",
x"009D",
x"0093",
x"008E",
x"0088",
x"007C",
x"0087",
x"008E",
x"0092",
x"009A",
x"0098",
x"00A0",
x"009B",
x"009E",
x"0052",
x"0024",
x"0017",
x"000F",
x"0005",
x"0007",
x"002F",
x"006C",
x"0099",
x"009C",
x"0092",
x"0095",
x"0087",
x"008C",
x"008F",
x"0081",
x"0081",
x"0086",
x"0092",
x"008B",
x"007D",
x"008F",
x"0095",
x"008C",
x"008B",
x"0000",
x"0000",
x"0000",
x"0000",
x"00B6",
x"00B7",
x"00B6",
x"00B5",
x"00B6",
x"00B7",
x"00B8",
x"00B5",
x"00B6",
x"00B6",
x"00B5",
x"00B7",
x"00B6",
x"00B6",
x"00B9",
x"00B8",
x"00B9",
x"00BA",
x"00B9",
x"00B8",
x"00B7",
x"00B8",
x"00B9",
x"00B7",
x"00B8",
x"00B9",
x"00B7",
x"00B7",
x"00B7",
x"00B5",
x"00B7",
x"00B8",
x"00B6",
x"00B6",
x"00B7",
x"00B7",
x"00B7",
x"00B8",
x"00B6",
x"00B5",
x"00B6",
x"00B5",
x"00B3",
x"00B4",
x"00B4",
x"00B4",
x"00B2",
x"00B3",
x"00B2",
x"00B1",
x"00B1",
x"00B2",
x"00B1",
x"00B1",
x"00B1",
x"00AF",
x"00B0",
x"00AF",
x"00AE",
x"00AE",
x"00B0",
x"00AF",
x"00AE",
x"00B0",
x"00B0",
x"00B0",
x"00AF",
x"00AE",
x"00AC",
x"00AE",
x"00B5",
x"00A7",
x"00AD",
x"00A7",
x"00A2",
x"00AD",
x"00C0",
x"00AF",
x"0096",
x"00B7",
x"00CC",
x"00B1",
x"004C",
x"0027",
x"0039",
x"0044",
x"0052",
x"0073",
x"0093",
x"00A0",
x"00A3",
x"0098",
x"008B",
x"0087",
x"007C",
x"0088",
x"008D",
x"008E",
x"0096",
x"0097",
x"009C",
x"009A",
x"0096",
x"009E",
x"0084",
x"0054",
x"002C",
x"001C",
x"0013",
x"0007",
x"0007",
x"0027",
x"0057",
x"0083",
x"0091",
x"008F",
x"0096",
x"008E",
x"0086",
x"0080",
x"008F",
x"008F",
x"008F",
x"0089",
x"0085",
x"008C",
x"0091",
x"0089",
x"0000",
x"0000",
x"0000",
x"0000",
x"00B7",
x"00B8",
x"00B7",
x"00B7",
x"00B6",
x"00B7",
x"00B8",
x"00B5",
x"00B6",
x"00B7",
x"00B4",
x"00B5",
x"00B6",
x"00B6",
x"00B8",
x"00B9",
x"00B9",
x"00B9",
x"00B8",
x"00B7",
x"00B6",
x"00B8",
x"00BA",
x"00B7",
x"00B7",
x"00B8",
x"00B7",
x"00B7",
x"00B6",
x"00B5",
x"00B6",
x"00B8",
x"00B6",
x"00B5",
x"00B7",
x"00B7",
x"00B7",
x"00B8",
x"00B5",
x"00B5",
x"00B6",
x"00B4",
x"00B2",
x"00B4",
x"00B4",
x"00B3",
x"00B2",
x"00B2",
x"00B2",
x"00B2",
x"00B2",
x"00B0",
x"00AF",
x"00B1",
x"00AF",
x"00AF",
x"00B0",
x"00AE",
x"00AF",
x"00AD",
x"00AF",
x"00AE",
x"00AF",
x"00B0",
x"00B0",
x"00AF",
x"00AF",
x"00AE",
x"00AD",
x"00AF",
x"00AF",
x"00AF",
x"00AF",
x"00AE",
x"00AD",
x"00AB",
x"00B9",
x"00B6",
x"00A3",
x"00B5",
x"00BB",
x"005F",
x"001B",
x"0024",
x"0028",
x"0031",
x"0057",
x"0079",
x"0094",
x"00A1",
x"009E",
x"0095",
x"0086",
x"0085",
x"007E",
x"008B",
x"008E",
x"008E",
x"0092",
x"009B",
x"009E",
x"009B",
x"0096",
x"0098",
x"009C",
x"0090",
x"007C",
x"005C",
x"0039",
x"001D",
x"0012",
x"000A",
x"0001",
x"003B",
x"0073",
x"006C",
x"0091",
x"0094",
x"0085",
x"0092",
x"0098",
x"008C",
x"0087",
x"008B",
x"0085",
x"008F",
x"008B",
x"007A",
x"0000",
x"0000",
x"0000",
x"0000",
x"00B7",
x"00B7",
x"00B5",
x"00B7",
x"00B6",
x"00B6",
x"00B7",
x"00B4",
x"00B7",
x"00B8",
x"00B5",
x"00B5",
x"00B6",
x"00B5",
x"00B6",
x"00B8",
x"00B8",
x"00B8",
x"00B7",
x"00B5",
x"00B6",
x"00B8",
x"00B9",
x"00B8",
x"00B8",
x"00B8",
x"00B6",
x"00B6",
x"00B6",
x"00B5",
x"00B6",
x"00B7",
x"00B6",
x"00B7",
x"00B9",
x"00B7",
x"00B4",
x"00B6",
x"00B5",
x"00B5",
x"00B6",
x"00B5",
x"00B3",
x"00B4",
x"00B6",
x"00B3",
x"00B2",
x"00B3",
x"00B2",
x"00B2",
x"00B1",
x"00AF",
x"00AF",
x"00AF",
x"00AF",
x"00B0",
x"00B1",
x"00AB",
x"00A5",
x"00A5",
x"00A6",
x"00A4",
x"00A5",
x"00A7",
x"00A4",
x"00A4",
x"00A6",
x"00A4",
x"00A4",
x"00A5",
x"00A4",
x"00A3",
x"00A4",
x"00A2",
x"00A1",
x"009F",
x"00AD",
x"00B7",
x"00A5",
x"009B",
x"0081",
x"002E",
x"001C",
x"0022",
x"002A",
x"0028",
x"0052",
x"007F",
x"0096",
x"00A3",
x"009E",
x"0093",
x"0088",
x"0084",
x"007B",
x"0087",
x"0091",
x"0094",
x"0095",
x"0092",
x"009C",
x"009B",
x"009A",
x"009A",
x"009B",
x"008B",
x"008F",
x"0090",
x"0090",
x"0074",
x"0043",
x"0025",
x"0019",
x"0093",
x"00C0",
x"0079",
x"0056",
x"0073",
x"0079",
x"0088",
x"008E",
x"0083",
x"007E",
x"008A",
x"0088",
x"007E",
x"008E",
x"0081",
x"0000",
x"0000",
x"0000",
x"0000",
x"00B6",
x"00B6",
x"00B6",
x"00B7",
x"00B7",
x"00B8",
x"00B7",
x"00B7",
x"00B6",
x"00B6",
x"00B6",
x"00B5",
x"00B5",
x"00B3",
x"00B7",
x"00B8",
x"00B8",
x"00B8",
x"00B6",
x"00B6",
x"00B8",
x"00B8",
x"00B9",
x"00B8",
x"00B7",
x"00BA",
x"00B6",
x"00B6",
x"00B6",
x"00B5",
x"00B6",
x"00B6",
x"00B6",
x"00B6",
x"00B9",
x"00B6",
x"00B4",
x"00B6",
x"00B5",
x"00B5",
x"00B6",
x"00B4",
x"00B2",
x"00B4",
x"00B5",
x"00B4",
x"00B2",
x"00B4",
x"00B4",
x"00B1",
x"00B0",
x"00AE",
x"00AF",
x"00AE",
x"00B0",
x"00A6",
x"0092",
x"00B2",
x"00BE",
x"00BE",
x"00BC",
x"00BA",
x"00BA",
x"00BB",
x"00B9",
x"00B9",
x"00B9",
x"00B8",
x"00B9",
x"00B8",
x"00B7",
x"00B5",
x"00B2",
x"00B1",
x"00B4",
x"00B2",
x"00B6",
x"00AF",
x"0084",
x"0080",
x"0078",
x"002A",
x"0021",
x"0026",
x"0030",
x"0033",
x"005A",
x"0079",
x"0097",
x"00A4",
x"009F",
x"0098",
x"0087",
x"007E",
x"007B",
x"0087",
x"0090",
x"0091",
x"0093",
x"0094",
x"009C",
x"0095",
x"0099",
x"0098",
x"0098",
x"008F",
x"008D",
x"008B",
x"0094",
x"00A5",
x"0091",
x"0071",
x"006B",
x"00E2",
x"00E7",
x"00B0",
x"006A",
x"0049",
x"0046",
x"0062",
x"0094",
x"0098",
x"008D",
x"00A5",
x"0092",
x"008A",
x"008D",
x"0077",
x"0000",
x"0000",
x"0000",
x"0000",
x"00B5",
x"00B5",
x"00B6",
x"00B7",
x"00B7",
x"00B8",
x"00B7",
x"00B5",
x"00B8",
x"00B7",
x"00B6",
x"00B7",
x"00B7",
x"00B7",
x"00B7",
x"00B8",
x"00B6",
x"00B7",
x"00B8",
x"00B7",
x"00B6",
x"00B7",
x"00B7",
x"00B7",
x"00B8",
x"00B8",
x"00B4",
x"00B6",
x"00B7",
x"00B5",
x"00B6",
x"00B7",
x"00B6",
x"00B5",
x"00B6",
x"00B6",
x"00B5",
x"00B6",
x"00B4",
x"00B4",
x"00B7",
x"00B5",
x"00B3",
x"00B5",
x"00B4",
x"00B3",
x"00B3",
x"00B4",
x"00B4",
x"00B2",
x"00B1",
x"00B0",
x"00B0",
x"00B1",
x"00B3",
x"009F",
x"007A",
x"00B1",
x"00C8",
x"00C7",
x"00C8",
x"00C7",
x"00C8",
x"00C6",
x"00C4",
x"00C4",
x"00C4",
x"00C2",
x"00C4",
x"00C3",
x"00C1",
x"00C1",
x"00BF",
x"00BF",
x"00C5",
x"00C4",
x"00C1",
x"00A7",
x"0070",
x"008C",
x"0089",
x"0034",
x"0028",
x"002B",
x"002D",
x"0041",
x"0083",
x"008A",
x"0096",
x"00A4",
x"00A1",
x"0096",
x"0083",
x"007C",
x"0077",
x"0082",
x"008E",
x"0094",
x"0097",
x"0099",
x"009F",
x"0095",
x"0099",
x"0090",
x"008A",
x"008B",
x"0093",
x"008E",
x"0097",
x"00A3",
x"0088",
x"0097",
x"0098",
x"00AC",
x"00C5",
x"00AB",
x"00D6",
x"00C5",
x"0087",
x"0052",
x"004E",
x"0064",
x"0079",
x"0091",
x"0083",
x"008D",
x"0086",
x"008E",
x"0000",
x"0000",
x"0000",
x"0000",
x"00B5",
x"00B5",
x"00B6",
x"00B5",
x"00B6",
x"00B6",
x"00B7",
x"00B5",
x"00B8",
x"00B8",
x"00B5",
x"00B6",
x"00B5",
x"00B6",
x"00B7",
x"00B8",
x"00B6",
x"00B6",
x"00B8",
x"00B7",
x"00B6",
x"00B7",
x"00B8",
x"00B7",
x"00B8",
x"00B8",
x"00B5",
x"00B4",
x"00B5",
x"00B5",
x"00B4",
x"00B6",
x"00B6",
x"00B3",
x"00B4",
x"00B3",
x"00B3",
x"00B5",
x"00B4",
x"00B4",
x"00B4",
x"00B4",
x"00B3",
x"00B5",
x"00B3",
x"00B2",
x"00B2",
x"00B4",
x"00B4",
x"00B2",
x"00B2",
x"00AF",
x"00AD",
x"00AC",
x"00A6",
x"0097",
x"0087",
x"00B7",
x"00C6",
x"00C5",
x"00C6",
x"00C6",
x"00C7",
x"00C4",
x"00C4",
x"00C2",
x"00C0",
x"00BF",
x"00C0",
x"00C1",
x"00C0",
x"00BF",
x"00BF",
x"00BE",
x"00BF",
x"00BE",
x"00BD",
x"00AC",
x"0089",
x"00A2",
x"009D",
x"0041",
x"002A",
x"0031",
x"0030",
x"0031",
x"006C",
x"008A",
x"0098",
x"00A6",
x"00A1",
x"0098",
x"0085",
x"007B",
x"007A",
x"007E",
x"008F",
x"0092",
x"0095",
x"0096",
x"009E",
x"0099",
x"0097",
x"0086",
x"0083",
x"008C",
x"0093",
x"008B",
x"0096",
x"009C",
x"008F",
x"0090",
x"0093",
x"0092",
x"009C",
x"0084",
x"0099",
x"00B5",
x"00D5",
x"00D1",
x"009B",
x"005E",
x"004A",
x"0059",
x"0078",
x"0091",
x"008F",
x"008A",
x"0000",
x"0000",
x"0000",
x"0000",
x"00B5",
x"00B5",
x"00B6",
x"00B3",
x"00B3",
x"00B6",
x"00B6",
x"00B5",
x"00B6",
x"00B7",
x"00B6",
x"00B5",
x"00B7",
x"00B6",
x"00B6",
x"00B7",
x"00B5",
x"00B5",
x"00B7",
x"00B6",
x"00B4",
x"00B7",
x"00B6",
x"00B4",
x"00B7",
x"00B7",
x"00B5",
x"00B5",
x"00B4",
x"00B3",
x"00B3",
x"00B4",
x"00B3",
x"00B3",
x"00B3",
x"00B1",
x"00B1",
x"00B3",
x"00B3",
x"00B2",
x"00B3",
x"00B4",
x"00B2",
x"00B3",
x"00B3",
x"00B2",
x"00B2",
x"00B3",
x"00B1",
x"00AF",
x"00B2",
x"00B0",
x"00AC",
x"00B2",
x"00BF",
x"009C",
x"0072",
x"00B0",
x"00C7",
x"00C6",
x"00C4",
x"00C6",
x"00C4",
x"00C4",
x"00C4",
x"00C3",
x"00C1",
x"00BE",
x"00C0",
x"00C2",
x"00C2",
x"00C0",
x"00C1",
x"00BF",
x"00BA",
x"00BD",
x"00BE",
x"00B1",
x"0094",
x"00AA",
x"00B1",
x"005D",
x"002A",
x"0035",
x"0046",
x"0035",
x"0054",
x"007C",
x"009A",
x"00A4",
x"00A1",
x"0095",
x"0087",
x"007A",
x"0077",
x"007D",
x"008D",
x"008B",
x"0093",
x"0092",
x"0094",
x"0090",
x"0096",
x"0097",
x"008B",
x"0085",
x"0090",
x"008A",
x"008B",
x"0096",
x"008E",
x"0086",
x"008E",
x"0091",
x"0091",
x"008A",
x"008C",
x"0077",
x"008C",
x"00AC",
x"00C9",
x"00D5",
x"00B4",
x"0073",
x"0050",
x"0059",
x"007A",
x"0094",
x"0000",
x"0000",
x"0000",
x"0000",
x"00B6",
x"00B7",
x"00B6",
x"00B3",
x"00B3",
x"00B6",
x"00B5",
x"00B3",
x"00B6",
x"00B6",
x"00B4",
x"00B5",
x"00B6",
x"00B4",
x"00B5",
x"00B6",
x"00B5",
x"00B6",
x"00B7",
x"00B5",
x"00B5",
x"00B7",
x"00B5",
x"00B4",
x"00B6",
x"00B6",
x"00B4",
x"00B4",
x"00B4",
x"00B3",
x"00B3",
x"00B4",
x"00B2",
x"00B3",
x"00B3",
x"00B1",
x"00B0",
x"00B2",
x"00B2",
x"00B2",
x"00B3",
x"00B3",
x"00B2",
x"00B3",
x"00B4",
x"00B1",
x"00B2",
x"00B2",
x"00B1",
x"00B1",
x"00B2",
x"00B0",
x"00AE",
x"00BD",
x"00DD",
x"00C1",
x"0097",
x"00B9",
x"00C5",
x"00C4",
x"00C6",
x"00C7",
x"00C5",
x"00C5",
x"00C4",
x"00C5",
x"00C5",
x"00C1",
x"00C4",
x"00C6",
x"00C5",
x"00C4",
x"00C4",
x"00C3",
x"00C3",
x"00C4",
x"00C1",
x"00B3",
x"009D",
x"00AC",
x"00BE",
x"0085",
x"002F",
x"0038",
x"003F",
x"0036",
x"005A",
x"007E",
x"0099",
x"00A2",
x"00A2",
x"0094",
x"0084",
x"0077",
x"0074",
x"0080",
x"008D",
x"008F",
x"008E",
x"0095",
x"0093",
x"0090",
x"0099",
x"009E",
x"008C",
x"007B",
x"0090",
x"008C",
x"0093",
x"0094",
x"0096",
x"0087",
x"0088",
x"0090",
x"0090",
x"008A",
x"008A",
x"007B",
x"008B",
x"008B",
x"008C",
x"009E",
x"00C7",
x"00DC",
x"00BB",
x"007D",
x"004F",
x"004C",
x"0000",
x"0000",
x"0000",
x"0000",
x"00B6",
x"00B6",
x"00B6",
x"00B5",
x"00B3",
x"00B4",
x"00B6",
x"00B3",
x"00B4",
x"00B4",
x"00B3",
x"00B5",
x"00B6",
x"00B5",
x"00B5",
x"00B6",
x"00B5",
x"00B5",
x"00B6",
x"00B3",
x"00B5",
x"00B6",
x"00B5",
x"00B4",
x"00B6",
x"00B6",
x"00B4",
x"00B5",
x"00B4",
x"00B3",
x"00B2",
x"00B4",
x"00B1",
x"00B2",
x"00B2",
x"00B1",
x"00B2",
x"00B3",
x"00B3",
x"00B3",
x"00B3",
x"00B2",
x"00B1",
x"00B2",
x"00B2",
x"00B1",
x"00B1",
x"00B2",
x"00B1",
x"00B1",
x"00B2",
x"00B1",
x"00AF",
x"00B3",
x"00C3",
x"00BC",
x"00AF",
x"00B9",
x"00C0",
x"00C1",
x"00C2",
x"00C4",
x"00C2",
x"00C2",
x"00C2",
x"00C2",
x"00C3",
x"00C1",
x"00C3",
x"00C5",
x"00C4",
x"00C4",
x"00C5",
x"00C5",
x"00C8",
x"00C7",
x"00C1",
x"00B1",
x"00A4",
x"00B0",
x"00C0",
x"00B1",
x"0044",
x"002F",
x"0034",
x"0031",
x"004B",
x"007E",
x"009B",
x"00A3",
x"00A2",
x"0094",
x"0089",
x"007E",
x"0075",
x"0084",
x"008F",
x"008E",
x"008F",
x"0096",
x"0095",
x"008D",
x"0092",
x"0098",
x"0090",
x"007F",
x"008A",
x"008B",
x"0093",
x"009E",
x"0094",
x"008C",
x"008C",
x"008D",
x"009A",
x"0089",
x"0095",
x"007C",
x"0078",
x"0084",
x"0090",
x"007B",
x"007F",
x"009D",
x"00B8",
x"00DA",
x"00C7",
x"0097",
x"0000",
x"0000",
x"0000",
x"0000",
x"00B5",
x"00B5",
x"00B6",
x"00B5",
x"00B4",
x"00B5",
x"00B4",
x"00B2",
x"00B5",
x"00B4",
x"00B3",
x"00B5",
x"00B5",
x"00B3",
x"00B5",
x"00B6",
x"00B4",
x"00B4",
x"00B4",
x"00B4",
x"00B4",
x"00B4",
x"00B4",
x"00B3",
x"00B5",
x"00B7",
x"00B3",
x"00B4",
x"00B3",
x"00B1",
x"00B2",
x"00B4",
x"00B1",
x"00B1",
x"00B2",
x"00B1",
x"00B1",
x"00B3",
x"00B3",
x"00B3",
x"00B3",
x"00B1",
x"00B0",
x"00B1",
x"00B2",
x"00B2",
x"00B1",
x"00B2",
x"00B3",
x"00B1",
x"00B0",
x"00AF",
x"00AE",
x"00AE",
x"00AD",
x"00AE",
x"00AE",
x"00AF",
x"00AF",
x"00AF",
x"00AF",
x"00B0",
x"00AE",
x"00B1",
x"00B0",
x"00B1",
x"00B1",
x"00AF",
x"00AF",
x"00AD",
x"00AF",
x"00B1",
x"00B1",
x"00B0",
x"00B2",
x"00B1",
x"00B4",
x"00B0",
x"00A7",
x"00B4",
x"00C3",
x"00C8",
x"0071",
x"0026",
x"002D",
x"002B",
x"0044",
x"007B",
x"009D",
x"00A4",
x"00A3",
x"0099",
x"0088",
x"0079",
x"0071",
x"007F",
x"008A",
x"0087",
x"0091",
x"0094",
x"0097",
x"008C",
x"0090",
x"008D",
x"008B",
x"007B",
x"0087",
x"007E",
x"0080",
x"0099",
x"008A",
x"008E",
x"008F",
x"0088",
x"0090",
x"007F",
x"008C",
x"008F",
x"0084",
x"0083",
x"0088",
x"0086",
x"0089",
x"0090",
x"007F",
x"008B",
x"00AC",
x"00D0",
x"0000",
x"0000",
x"0000",
x"0000",
x"00B6",
x"00B6",
x"00B6",
x"00B5",
x"00B5",
x"00B4",
x"00B5",
x"00B3",
x"00B4",
x"00B5",
x"00B2",
x"00B4",
x"00B4",
x"00B3",
x"00B4",
x"00B5",
x"00B3",
x"00B3",
x"00B4",
x"00B4",
x"00B3",
x"00B4",
x"00B3",
x"00B2",
x"00B4",
x"00B5",
x"00B2",
x"00B1",
x"00B2",
x"00B1",
x"00B1",
x"00B2",
x"00B1",
x"00B1",
x"00B2",
x"00B1",
x"00B1",
x"00B3",
x"00B2",
x"00B1",
x"00B3",
x"00B1",
x"00B0",
x"00B4",
x"00B3",
x"00B1",
x"00B1",
x"00B1",
x"00B1",
x"00B0",
x"00AF",
x"00AF",
x"00AF",
x"00B0",
x"00AF",
x"00AD",
x"00AE",
x"00AE",
x"00AE",
x"00AE",
x"00AF",
x"00AE",
x"00AF",
x"00AE",
x"00AE",
x"00B0",
x"00AE",
x"00AD",
x"00AD",
x"00AC",
x"00AC",
x"00AE",
x"00AE",
x"00AB",
x"00AB",
x"00AC",
x"00AD",
x"00A8",
x"00AA",
x"00BC",
x"00C4",
x"00C9",
x"00A7",
x"0035",
x"0025",
x"002C",
x"004D",
x"0083",
x"009D",
x"00A3",
x"00A3",
x"0099",
x"0088",
x"0075",
x"0075",
x"0081",
x"0088",
x"008D",
x"0090",
x"008E",
x"0097",
x"008C",
x"0088",
x"0089",
x"0089",
x"0086",
x"008D",
x"0087",
x"0081",
x"008B",
x"007C",
x"008B",
x"008E",
x"0088",
x"008E",
x"0080",
x"0088",
x"0088",
x"008D",
x"008E",
x"0086",
x"0088",
x"008A",
x"0091",
x"0086",
x"0081",
x"0080",
x"00A0",
x"0000",
x"0000",
x"0000",
x"0000",
x"00B6",
x"00B6",
x"00B5",
x"00B5",
x"00B5",
x"00B6",
x"00B4",
x"00B3",
x"00B5",
x"00B4",
x"00B3",
x"00B3",
x"00B4",
x"00B4",
x"00B3",
x"00B4",
x"00B3",
x"00B3",
x"00B5",
x"00B2",
x"00B1",
x"00B3",
x"00B3",
x"00B3",
x"00B4",
x"00B2",
x"00B0",
x"00B2",
x"00B1",
x"00B0",
x"00B0",
x"00B1",
x"00B0",
x"00B2",
x"00B1",
x"00AF",
x"00B0",
x"00B1",
x"00B2",
x"00B1",
x"00B2",
x"00B1",
x"00B0",
x"00B0",
x"00B2",
x"00B1",
x"00B2",
x"00B1",
x"00B1",
x"00B0",
x"00AE",
x"00AE",
x"00AE",
x"00AE",
x"00AF",
x"00AD",
x"00AF",
x"00AE",
x"00AE",
x"00AE",
x"00AF",
x"00AD",
x"00B0",
x"00AF",
x"00AF",
x"00AF",
x"00AF",
x"00AC",
x"00AC",
x"00AC",
x"00AC",
x"00AD",
x"00AD",
x"00AC",
x"00AB",
x"00AB",
x"00AD",
x"00A8",
x"00B1",
x"00C1",
x"00C3",
x"00C8",
x"00C6",
x"0071",
x"0025",
x"0030",
x"0058",
x"0085",
x"009C",
x"009F",
x"009F",
x"0095",
x"0084",
x"0078",
x"0078",
x"007F",
x"0088",
x"0092",
x"0091",
x"008D",
x"0093",
x"008D",
x"008D",
x"008C",
x"008D",
x"007F",
x"008C",
x"0081",
x"007B",
x"008D",
x"0088",
x"007F",
x"008F",
x"0091",
x"008E",
x"0078",
x"007B",
x"0080",
x"008A",
x"007E",
x"0087",
x"008E",
x"0091",
x"008C",
x"0090",
x"0086",
x"006F",
x"0098",
x"0000",
x"0000",
x"0000",
x"0000",
x"00B4",
x"00B4",
x"00B4",
x"00B2",
x"00B3",
x"00B6",
x"00B5",
x"00B3",
x"00B5",
x"00B5",
x"00B2",
x"00B3",
x"00B1",
x"00B0",
x"00B2",
x"00B3",
x"00B1",
x"00B2",
x"00B5",
x"00B3",
x"00B1",
x"00B2",
x"00B1",
x"00B2",
x"00B2",
x"00B2",
x"00B1",
x"00B1",
x"00B0",
x"00AE",
x"00B1",
x"00B1",
x"00B1",
x"00B2",
x"00B1",
x"00AF",
x"00AF",
x"00B1",
x"00B0",
x"00B1",
x"00B2",
x"00B1",
x"00B0",
x"00B2",
x"00B1",
x"00B0",
x"00B1",
x"00B2",
x"00B1",
x"00AF",
x"00AE",
x"00AD",
x"00AF",
x"00B1",
x"00AD",
x"00AC",
x"00AF",
x"00AE",
x"00AD",
x"00AF",
x"00AF",
x"00B0",
x"00AF",
x"00AF",
x"00AE",
x"00AE",
x"00AD",
x"00AC",
x"00AC",
x"00AD",
x"00AC",
x"00AB",
x"00AC",
x"00AC",
x"00AA",
x"00AA",
x"00A9",
x"00A9",
x"00B8",
x"00C1",
x"00C1",
x"00C8",
x"00CB",
x"00B3",
x"0045",
x"0027",
x"0062",
x"0085",
x"009C",
x"009F",
x"00A1",
x"0095",
x"0081",
x"0077",
x"0077",
x"007D",
x"0082",
x"008D",
x"0092",
x"0091",
x"0093",
x"008D",
x"0093",
x"0091",
x"0090",
x"0088",
x"0082",
x"008B",
x"0083",
x"0092",
x"008A",
x"007E",
x"0084",
x"008B",
x"008C",
x"0080",
x"0095",
x"0087",
x"0082",
x"0080",
x"0086",
x"0083",
x"008F",
x"0097",
x"0091",
x"008C",
x"0072",
x"007C",
x"0000",
x"0000",
x"0000",
x"0000",
x"00B3",
x"00B3",
x"00B3",
x"00B1",
x"00B1",
x"00B4",
x"00B4",
x"00B2",
x"00B5",
x"00B4",
x"00B4",
x"00B3",
x"00B1",
x"00B1",
x"00B2",
x"00B2",
x"00B2",
x"00B2",
x"00B3",
x"00B2",
x"00B1",
x"00B2",
x"00B1",
x"00B2",
x"00B2",
x"00B1",
x"00B1",
x"00B1",
x"00B2",
x"00AE",
x"00AF",
x"00B0",
x"00AF",
x"00AF",
x"00B1",
x"00AF",
x"00B0",
x"00B1",
x"00B0",
x"00B0",
x"00B1",
x"00B0",
x"00B0",
x"00B1",
x"00B1",
x"00AF",
x"00B1",
x"00B0",
x"00B0",
x"00AF",
x"00AF",
x"00AE",
x"00AE",
x"00AE",
x"00AD",
x"00AD",
x"00AD",
x"00AE",
x"00AF",
x"00B0",
x"00AE",
x"00AF",
x"00B0",
x"00B0",
x"00AE",
x"00AF",
x"00AF",
x"00AC",
x"00AD",
x"00AE",
x"00AC",
x"00AD",
x"00AD",
x"00AB",
x"00AC",
x"00AC",
x"00A5",
x"00A8",
x"00B9",
x"00C4",
x"00C5",
x"00C8",
x"00CD",
x"00CB",
x"008F",
x"0032",
x"006E",
x"008B",
x"009C",
x"009F",
x"009F",
x"0096",
x"0083",
x"0075",
x"0078",
x"0080",
x"008B",
x"008D",
x"0092",
x"0095",
x"0095",
x"008A",
x"008B",
x"008D",
x"0090",
x"0088",
x"0080",
x"008A",
x"008D",
x"008F",
x"0084",
x"0091",
x"0084",
x"007E",
x"0087",
x"008A",
x"0091",
x"0076",
x"0085",
x"007C",
x"0072",
x"0080",
x"0096",
x"009B",
x"0090",
x"0092",
x"0078",
x"0063",
x"0000",
x"0000",
x"0000",
x"0000",
x"00B2",
x"00B2",
x"00B1",
x"00B0",
x"00B0",
x"00B4",
x"00B4",
x"00B2",
x"00B2",
x"00B3",
x"00B2",
x"00B1",
x"00B2",
x"00B1",
x"00B2",
x"00B1",
x"00B0",
x"00B0",
x"00B2",
x"00B1",
x"00B0",
x"00B1",
x"00B1",
x"00B1",
x"00B1",
x"00B0",
x"00B1",
x"00B1",
x"00B0",
x"00B0",
x"00AF",
x"00B1",
x"00AF",
x"00AE",
x"00AF",
x"00B0",
x"00AF",
x"00B0",
x"00AF",
x"00AE",
x"00AF",
x"00AD",
x"00AC",
x"00B0",
x"00AF",
x"00AD",
x"00B1",
x"00B0",
x"00AD",
x"00AD",
x"00AE",
x"00AE",
x"00AE",
x"00AE",
x"00AE",
x"00AD",
x"00AD",
x"00AD",
x"00AF",
x"00AE",
x"00AE",
x"00AE",
x"00AF",
x"00AF",
x"00AD",
x"00AE",
x"00AD",
x"00AC",
x"00AC",
x"00AD",
x"00AC",
x"00AE",
x"00AE",
x"00AB",
x"00AB",
x"00AD",
x"00A1",
x"00A7",
x"00B9",
x"00C2",
x"00C3",
x"00C7",
x"00CC",
x"00C5",
x"00BB",
x"006B",
x"0062",
x"008C",
x"009D",
x"00A0",
x"009F",
x"0094",
x"0083",
x"0074",
x"0079",
x"007A",
x"008D",
x"008D",
x"008F",
x"0092",
x"008E",
x"008F",
x"008E",
x"0085",
x"008B",
x"008C",
x"0091",
x"0090",
x"008F",
x"008B",
x"0088",
x"007E",
x"0088",
x"008B",
x"008B",
x"007B",
x"008E",
x"0077",
x"0077",
x"0088",
x"0079",
x"007C",
x"008F",
x"0094",
x"008E",
x"008E",
x"0078",
x"0078",
x"0000",
x"0000",
x"0000",
x"0000",
x"00B2",
x"00B2",
x"00B0",
x"00AF",
x"00B0",
x"00B2",
x"00B3",
x"00B1",
x"00B2",
x"00B3",
x"00B0",
x"00B1",
x"00B0",
x"00AE",
x"00B0",
x"00B0",
x"00B0",
x"00B1",
x"00B1",
x"00B0",
x"00AF",
x"00B0",
x"00B0",
x"00B1",
x"00B0",
x"00B1",
x"00AF",
x"00B0",
x"00B0",
x"00AF",
x"00AF",
x"00AE",
x"00AD",
x"00AD",
x"00AD",
x"00AD",
x"00AD",
x"00AE",
x"00AE",
x"00AD",
x"00AE",
x"00AF",
x"00AB",
x"00AE",
x"00AE",
x"00AC",
x"00AE",
x"00AE",
x"00AD",
x"00AD",
x"00AD",
x"00AC",
x"00AC",
x"00AD",
x"00AB",
x"00AB",
x"00AC",
x"00AD",
x"00AE",
x"00AE",
x"00AE",
x"00AD",
x"00AE",
x"00AD",
x"00AD",
x"00AC",
x"00AC",
x"00AB",
x"00AB",
x"00AE",
x"00AD",
x"00AD",
x"00AD",
x"00AD",
x"00AD",
x"00AD",
x"00A0",
x"00A9",
x"00BB",
x"00C4",
x"00C5",
x"00C6",
x"00CC",
x"00C7",
x"00C1",
x"0091",
x"0071",
x"008A",
x"009C",
x"009F",
x"00A0",
x"0094",
x"007C",
x"0071",
x"007A",
x"007A",
x"0090",
x"0092",
x"008A",
x"0095",
x"0092",
x"008A",
x"0088",
x"0080",
x"0085",
x"008C",
x"008C",
x"0093",
x"0086",
x"008B",
x"008F",
x"0088",
x"008C",
x"008E",
x"0093",
x"007B",
x"0080",
x"007B",
x"0088",
x"0098",
x"0092",
x"0081",
x"0082",
x"008D",
x"009B",
x"0094",
x"0088",
x"0081",
x"0000",
x"0000",
x"0000",
x"0000",
x"00B0",
x"00B0",
x"00B1",
x"00AF",
x"00AD",
x"00AF",
x"00B1",
x"00B1",
x"00B2",
x"00B2",
x"00B0",
x"00B0",
x"00B0",
x"00AE",
x"00AF",
x"00B0",
x"00AE",
x"00B0",
x"00B0",
x"00AF",
x"00AE",
x"00B0",
x"00B0",
x"00AE",
x"00AF",
x"00AF",
x"00AE",
x"00B0",
x"00AF",
x"00AB",
x"00AC",
x"00AC",
x"00AC",
x"00AD",
x"00AC",
x"00AC",
x"00AB",
x"00AC",
x"00AD",
x"00AD",
x"00AD",
x"00AD",
x"00AA",
x"00AD",
x"00AD",
x"00AB",
x"00AC",
x"00AD",
x"00AB",
x"00AC",
x"00AC",
x"00AA",
x"00AB",
x"00AC",
x"00AA",
x"00AB",
x"00AC",
x"00AE",
x"00AE",
x"00AD",
x"00AE",
x"00AD",
x"00AD",
x"00AC",
x"00AC",
x"00AC",
x"00AC",
x"00B9",
x"00B0",
x"00AC",
x"00AE",
x"00AC",
x"00AD",
x"00AB",
x"00AB",
x"00AD",
x"00A2",
x"00AA",
x"00BA",
x"00C2",
x"00C6",
x"00C6",
x"00CD",
x"00CA",
x"00AC",
x"0071",
x"0073",
x"0085",
x"009B",
x"009F",
x"009F",
x"0093",
x"007B",
x"0070",
x"007D",
x"007C",
x"008F",
x"0092",
x"0089",
x"008E",
x"0090",
x"0089",
x"0088",
x"0089",
x"008B",
x"008B",
x"0080",
x"008C",
x"007F",
x"008C",
x"0091",
x"0094",
x"0091",
x"008B",
x"0095",
x"007E",
x"0084",
x"0079",
x"007D",
x"0082",
x"008A",
x"0090",
x"007F",
x"0091",
x"009C",
x"008D",
x"007C",
x"007E",
x"0000",
x"0000",
x"0000",
x"0000",
x"00B0",
x"00B1",
x"00B2",
x"00AF",
x"00AD",
x"00AE",
x"00B0",
x"00AF",
x"00B1",
x"00B1",
x"00AF",
x"00B0",
x"00B0",
x"00AE",
x"00B0",
x"00AE",
x"00AD",
x"00B0",
x"00B1",
x"00AC",
x"00AE",
x"00AF",
x"00AF",
x"00AD",
x"00AE",
x"00AE",
x"00AE",
x"00AF",
x"00AD",
x"00AC",
x"00AD",
x"00AC",
x"00AC",
x"00AE",
x"00AD",
x"00AB",
x"00AC",
x"00AD",
x"00AB",
x"00AC",
x"00AC",
x"00AB",
x"00A9",
x"00AB",
x"00AC",
x"00AB",
x"00AB",
x"00AD",
x"00AC",
x"00AB",
x"00AC",
x"00AA",
x"00AB",
x"00AB",
x"00AB",
x"00AB",
x"00AB",
x"00AC",
x"00AD",
x"00AD",
x"00AD",
x"00AD",
x"00AC",
x"00AB",
x"00AB",
x"00AA",
x"00B7",
x"00CB",
x"00B7",
x"00A3",
x"00A7",
x"00A7",
x"00A7",
x"00A4",
x"00A2",
x"00A1",
x"00A3",
x"00B0",
x"00BC",
x"00C3",
x"00C5",
x"00C7",
x"00CC",
x"00BE",
x"0071",
x"0057",
x"0082",
x"008B",
x"009B",
x"009F",
x"009E",
x"008F",
x"0077",
x"006F",
x"007D",
x"007C",
x"008F",
x"008E",
x"0090",
x"0092",
x"008D",
x"0084",
x"008D",
x"0087",
x"0088",
x"008D",
x"0079",
x"0089",
x"008A",
x"0091",
x"008A",
x"0085",
x"0090",
x"0091",
x"0094",
x"0075",
x"0078",
x"0076",
x"0073",
x"008D",
x"008A",
x"0093",
x"0090",
x"008A",
x"009B",
x"009A",
x"0082",
x"008A",
x"0000",
x"0000",
x"0000",
x"0000",
x"00B1",
x"00B1",
x"00B0",
x"00AE",
x"00AE",
x"00AF",
x"00B0",
x"00B0",
x"00B0",
x"00B1",
x"00AF",
x"00AF",
x"00AF",
x"00AE",
x"00B0",
x"00AD",
x"00AC",
x"00AE",
x"00B0",
x"00AC",
x"00AD",
x"00AF",
x"00AD",
x"00AD",
x"00AD",
x"00AE",
x"00AE",
x"00AD",
x"00AD",
x"00A9",
x"00AB",
x"00AC",
x"00AB",
x"00AC",
x"00AC",
x"00AB",
x"00AC",
x"00AB",
x"00AA",
x"00AB",
x"00AC",
x"00AA",
x"00AA",
x"00AB",
x"00AB",
x"00AA",
x"00AC",
x"00AC",
x"00AB",
x"00AB",
x"00AB",
x"00AA",
x"00AB",
x"00AA",
x"00AB",
x"00AA",
x"00AC",
x"00AB",
x"00AB",
x"00AC",
x"00AC",
x"00AB",
x"00AB",
x"00AB",
x"00A9",
x"00AC",
x"00C5",
x"00BE",
x"00AD",
x"00A8",
x"00A7",
x"00A6",
x"00A6",
x"00A5",
x"00A4",
x"00A4",
x"00A4",
x"00AD",
x"00BB",
x"00C2",
x"00C5",
x"00C8",
x"00C6",
x"008E",
x"004F",
x"005E",
x"006C",
x"0080",
x"009A",
x"009E",
x"009E",
x"008D",
x"0079",
x"006F",
x"007B",
x"007E",
x"008F",
x"008F",
x"008D",
x"0093",
x"008F",
x"0082",
x"0083",
x"007D",
x"0083",
x"008A",
x"007D",
x"0091",
x"0084",
x"0098",
x"0089",
x"0083",
x"008E",
x"0092",
x"008C",
x"0081",
x"0086",
x"0085",
x"0083",
x"008F",
x"0089",
x"008A",
x"0083",
x"008F",
x"0097",
x"008F",
x"007A",
x"008D",
x"0000",
x"0000",
x"0000",
x"0000",
x"00B0",
x"00B0",
x"00B0",
x"00AC",
x"00AC",
x"00AF",
x"00AF",
x"00B0",
x"00B1",
x"00B1",
x"00B0",
x"00B1",
x"00AE",
x"00AD",
x"00B0",
x"00AF",
x"00AC",
x"00AF",
x"00AF",
x"00AC",
x"00AC",
x"00AE",
x"00AC",
x"00AD",
x"00AD",
x"00AC",
x"00AC",
x"00AD",
x"00AC",
x"00A9",
x"00AA",
x"00AB",
x"00A7",
x"00A9",
x"00AA",
x"00A9",
x"00AB",
x"00AC",
x"00A9",
x"00AA",
x"00AB",
x"00AA",
x"00A9",
x"00AA",
x"00AA",
x"00A8",
x"00AB",
x"00AA",
x"00A9",
x"00AB",
x"00AA",
x"00A8",
x"00AA",
x"00A9",
x"00AA",
x"00AA",
x"00AC",
x"00AA",
x"00A9",
x"00A9",
x"00AB",
x"00AA",
x"00AB",
x"00AB",
x"00AA",
x"00AC",
x"00C2",
x"00C1",
x"00AD",
x"00A6",
x"00A4",
x"00A7",
x"00A4",
x"00A3",
x"00A3",
x"00A2",
x"00A5",
x"00B0",
x"00BC",
x"00C5",
x"00C6",
x"00CA",
x"00B2",
x"0055",
x"004E",
x"005E",
x"006D",
x"007B",
x"0098",
x"009D",
x"009D",
x"0091",
x"0078",
x"0071",
x"007A",
x"0080",
x"008D",
x"008A",
x"008D",
x"0093",
x"0093",
x"0085",
x"0084",
x"007E",
x"0089",
x"008D",
x"0078",
x"008E",
x"007F",
x"0093",
x"008F",
x"0087",
x"0088",
x"0087",
x"0095",
x"008F",
x"008B",
x"0081",
x"0086",
x"0093",
x"007C",
x"0080",
x"007A",
x"007E",
x"008E",
x"0083",
x"0073",
x"0084",
x"0000",
x"0000",
x"0000",
x"0000",
x"00AF",
x"00AF",
x"00AF",
x"00AE",
x"00AE",
x"00B0",
x"00B0",
x"00AF",
x"00B0",
x"00B1",
x"00AF",
x"00B0",
x"00AE",
x"00AD",
x"00AF",
x"00AE",
x"00AD",
x"00AF",
x"00AF",
x"00AA",
x"00AB",
x"00AD",
x"00AC",
x"00AC",
x"00AC",
x"00AA",
x"00AA",
x"00AC",
x"00AC",
x"00A9",
x"00A9",
x"00A9",
x"00A7",
x"00A9",
x"00AB",
x"00AA",
x"00AA",
x"00AA",
x"00AA",
x"00A9",
x"00AB",
x"00AA",
x"00A7",
x"00A8",
x"00A9",
x"00A9",
x"00A9",
x"00A8",
x"00A7",
x"00AA",
x"00AA",
x"00A9",
x"00AA",
x"00A9",
x"00A9",
x"00A9",
x"00AA",
x"00A9",
x"00A9",
x"00AA",
x"00AB",
x"00AA",
x"00AA",
x"00AB",
x"00AB",
x"00AA",
x"00B0",
x"00C9",
x"00B4",
x"009F",
x"009F",
x"00A5",
x"00A4",
x"00A3",
x"00A2",
x"00A1",
x"00A8",
x"00B1",
x"00BB",
x"00C7",
x"00C5",
x"00C3",
x"0083",
x"003F",
x"0038",
x"0045",
x"006A",
x"007D",
x"0098",
x"009B",
x"009D",
x"0090",
x"0078",
x"0074",
x"0077",
x"007D",
x"008D",
x"008B",
x"008E",
x"0094",
x"008C",
x"0082",
x"008D",
x"0087",
x"0089",
x"0082",
x"0083",
x"0096",
x"0083",
x"008F",
x"0089",
x"0080",
x"008E",
x"0088",
x"0090",
x"0081",
x"0088",
x"0080",
x"0085",
x"008B",
x"008C",
x"007E",
x"0073",
x"007B",
x"008C",
x"008C",
x"0080",
x"0083",
x"0000",
x"0000",
x"0000",
x"0000",
x"00AD",
x"00AD",
x"00AF",
x"00AC",
x"00AD",
x"00AF",
x"00AF",
x"00AE",
x"00B1",
x"00B1",
x"00AE",
x"00AF",
x"00AD",
x"00AC",
x"00AE",
x"00AF",
x"00AD",
x"00AE",
x"00AF",
x"00AA",
x"00AC",
x"00AE",
x"00AE",
x"00AD",
x"00AB",
x"00AB",
x"00A9",
x"00AC",
x"00AC",
x"00AA",
x"00AA",
x"00A9",
x"00A7",
x"00A8",
x"00A8",
x"00AA",
x"00AA",
x"00A8",
x"00A8",
x"00A9",
x"00AA",
x"00A9",
x"00A7",
x"00A9",
x"00AA",
x"00A8",
x"00A8",
x"00A8",
x"00AA",
x"00A9",
x"00A9",
x"00A9",
x"00A8",
x"00A8",
x"00A8",
x"00A8",
x"00AA",
x"00AA",
x"00A9",
x"00A8",
x"00A8",
x"00AA",
x"00AA",
x"00AA",
x"00AB",
x"00AA",
x"00AB",
x"00C5",
x"00B2",
x"00A3",
x"00A2",
x"00A3",
x"00A3",
x"00A5",
x"00A3",
x"00A5",
x"00AE",
x"00B1",
x"00BC",
x"00C5",
x"00C7",
x"00B3",
x"006E",
x"005F",
x"0057",
x"0059",
x"0076",
x"0080",
x"0097",
x"009A",
x"009B",
x"0093",
x"007B",
x"0075",
x"007A",
x"007E",
x"008D",
x"0088",
x"008A",
x"0096",
x"0091",
x"0080",
x"0089",
x"008D",
x"0091",
x"0085",
x"0082",
x"008E",
x"008B",
x"0094",
x"0085",
x"008C",
x"009D",
x"008C",
x"0084",
x"0086",
x"0084",
x"007A",
x"0076",
x"0079",
x"007E",
x"0081",
x"007B",
x"008D",
x"0090",
x"0091",
x"0083",
x"0085",
x"0000",
x"0000",
x"0000",
x"0000",
x"00AB",
x"00AB",
x"00AD",
x"00AD",
x"00AC",
x"00AD",
x"00AE",
x"00AD",
x"00B0",
x"00AF",
x"00AE",
x"00AF",
x"00AD",
x"00AC",
x"00AD",
x"00AD",
x"00AB",
x"00AD",
x"00AF",
x"00AB",
x"00AA",
x"00AE",
x"00AC",
x"00AB",
x"00AB",
x"00AA",
x"00AB",
x"00AB",
x"00AB",
x"00A8",
x"00A9",
x"00A8",
x"00A7",
x"00A8",
x"00A8",
x"00A9",
x"00A9",
x"00A9",
x"00A8",
x"00A9",
x"00A9",
x"00A8",
x"00A7",
x"00A8",
x"00A7",
x"00A7",
x"00A8",
x"00A8",
x"00A8",
x"00A7",
x"00A8",
x"00A9",
x"00A8",
x"00A8",
x"00A7",
x"00A8",
x"00A9",
x"00A8",
x"00A9",
x"00A9",
x"00A8",
x"00A7",
x"00A8",
x"00A8",
x"00A9",
x"00AB",
x"00AA",
x"00B8",
x"00B3",
x"00AF",
x"00AE",
x"00AD",
x"00AC",
x"00AB",
x"00AB",
x"00A4",
x"00A5",
x"00AA",
x"00BA",
x"00C6",
x"00C2",
x"009B",
x"0076",
x"007B",
x"007C",
x"0078",
x"0079",
x"007C",
x"0095",
x"009B",
x"009B",
x"0095",
x"007B",
x"0075",
x"007D",
x"007B",
x"008A",
x"0086",
x"008D",
x"0097",
x"008C",
x"0081",
x"0087",
x"0088",
x"008E",
x"0086",
x"007D",
x"0093",
x"008A",
x"0099",
x"0087",
x"0087",
x"008C",
x"008C",
x"008D",
x"0078",
x"0080",
x"007D",
x"0078",
x"0078",
x"0087",
x"0082",
x"007D",
x"008E",
x"0081",
x"007F",
x"0082",
x"007B",
x"0000",
x"0000",
x"0000",
x"0000",
x"00AB",
x"00AB",
x"00AD",
x"00AC",
x"00AB",
x"00AC",
x"00AA",
x"00AB",
x"00B0",
x"00AD",
x"00AB",
x"00AD",
x"00AE",
x"00AB",
x"00AC",
x"00AD",
x"00AB",
x"00AC",
x"00AD",
x"00AA",
x"00AA",
x"00AC",
x"00A9",
x"00A8",
x"00A9",
x"00A7",
x"00A7",
x"00A9",
x"00A9",
x"00A6",
x"00A7",
x"00A7",
x"00A5",
x"00A7",
x"00A7",
x"00A7",
x"00A8",
x"00A9",
x"00A6",
x"00A8",
x"00A7",
x"00A6",
x"00A6",
x"00A8",
x"00A7",
x"00A7",
x"00A6",
x"00A7",
x"00A6",
x"00A6",
x"00A7",
x"00A7",
x"00A6",
x"00A7",
x"00A7",
x"00A7",
x"00A8",
x"00A7",
x"00A7",
x"00A7",
x"00A7",
x"00A8",
x"00A8",
x"00A7",
x"00A9",
x"00A9",
x"00A7",
x"00A7",
x"00A9",
x"00A9",
x"00A8",
x"00AB",
x"00AA",
x"00A8",
x"00A7",
x"00A5",
x"00AD",
x"009F",
x"00B0",
x"00C0",
x"00B6",
x"0084",
x"0077",
x"007B",
x"007E",
x"0072",
x"0081",
x"0080",
x"0096",
x"009E",
x"009A",
x"0095",
x"0082",
x"007B",
x"007D",
x"007F",
x"0087",
x"0083",
x"0086",
x"0095",
x"0088",
x"007D",
x"0084",
x"007F",
x"0089",
x"0091",
x"0082",
x"0095",
x"0096",
x"008E",
x"0080",
x"007E",
x"0086",
x"009B",
x"008E",
x"0077",
x"0080",
x"0074",
x"0075",
x"007E",
x"0084",
x"0075",
x"0080",
x"0081",
x"007B",
x"0078",
x"007D",
x"008A",
x"0000",
x"0000",
x"0000",
x"0000",
x"00AC",
x"00AD",
x"00AC",
x"00AA",
x"00AC",
x"00AB",
x"00AA",
x"00AC",
x"00AD",
x"00AA",
x"00AA",
x"00AD",
x"00AC",
x"00AA",
x"00AB",
x"00AA",
x"00A8",
x"00AA",
x"00AC",
x"00A8",
x"00A9",
x"00A9",
x"00A7",
x"00A8",
x"00A7",
x"00A7",
x"00A6",
x"00A8",
x"00A9",
x"00A7",
x"00A7",
x"00A7",
x"00A4",
x"00A5",
x"00A7",
x"00A7",
x"00A6",
x"00A7",
x"00A6",
x"00A6",
x"00A7",
x"00A6",
x"00A5",
x"00A7",
x"00A6",
x"00A5",
x"00A6",
x"00A7",
x"00A5",
x"00A4",
x"00A6",
x"00A7",
x"00A6",
x"00A5",
x"00A5",
x"00A7",
x"00A8",
x"00A6",
x"00A6",
x"00A6",
x"00A6",
x"00A6",
x"00A8",
x"00A7",
x"00A8",
x"00A8",
x"00A7",
x"00A7",
x"00A7",
x"00A7",
x"00A7",
x"00A8",
x"00A7",
x"00A7",
x"00A7",
x"00A6",
x"00B2",
x"00A3",
x"00A5",
x"00BC",
x"00A5",
x"007A",
x"0077",
x"0077",
x"0076",
x"0076",
x"0072",
x"0079",
x"0098",
x"009C",
x"009A",
x"0092",
x"0082",
x"007F",
x"007E",
x"007E",
x"008E",
x"0086",
x"008A",
x"0097",
x"0089",
x"0080",
x"0084",
x"0087",
x"008E",
x"008F",
x"0081",
x"0084",
x"0092",
x"0091",
x"008B",
x"0083",
x"008F",
x"008D",
x"008F",
x"007A",
x"0081",
x"007B",
x"0076",
x"0072",
x"0075",
x"007F",
x"007A",
x"0089",
x"008E",
x"0092",
x"0091",
x"0089",
x"0000",
x"0000",
x"0000",
x"0000",
x"00AC",
x"00AC",
x"00AB",
x"00A9",
x"00A9",
x"00AA",
x"00AB",
x"00AD",
x"00B0",
x"00AB",
x"00AB",
x"00AD",
x"00AC",
x"00AA",
x"00AB",
x"00AA",
x"00A9",
x"00AA",
x"00A9",
x"00A9",
x"00A9",
x"00A7",
x"00A7",
x"00A7",
x"00A6",
x"00A6",
x"00A6",
x"00A8",
x"00A7",
x"00A5",
x"00A7",
x"00A6",
x"00A3",
x"00A5",
x"00A5",
x"00A6",
x"00A6",
x"00A6",
x"00A6",
x"00A7",
x"00A8",
x"00A6",
x"00A4",
x"00A7",
x"00A7",
x"00A4",
x"00A5",
x"00A6",
x"00A5",
x"00A4",
x"00A5",
x"00A5",
x"00A6",
x"00A5",
x"00A5",
x"00A6",
x"00A6",
x"00A6",
x"00A6",
x"00A6",
x"00A6",
x"00A5",
x"00A6",
x"00A8",
x"00A7",
x"00A8",
x"00A6",
x"00A6",
x"00A7",
x"00A7",
x"00A6",
x"00A7",
x"00A7",
x"00A7",
x"00A7",
x"00A5",
x"00AF",
x"00A1",
x"009F",
x"00B8",
x"0097",
x"0073",
x"0075",
x"0077",
x"0074",
x"006C",
x"004F",
x"0064",
x"0099",
x"009E",
x"009B",
x"0091",
x"0086",
x"0086",
x"0084",
x"0083",
x"008E",
x"0086",
x"0084",
x"0092",
x"0083",
x"0086",
x"0082",
x"0088",
x"0090",
x"008B",
x"007D",
x"007B",
x"008D",
x"009D",
x"0085",
x"007F",
x"0083",
x"0087",
x"008C",
x"0079",
x"0087",
x"0076",
x"007D",
x"0080",
x"0085",
x"0083",
x"007D",
x"0089",
x"0082",
x"0082",
x"0080",
x"0092",
x"0000",
x"0000",
x"0000",
x"0000",
x"00AA",
x"00AA",
x"00A9",
x"00A8",
x"00A7",
x"00A9",
x"00AB",
x"00AB",
x"00AD",
x"00AC",
x"00A9",
x"00AC",
x"00AA",
x"00AA",
x"00AB",
x"00AA",
x"00A8",
x"00A9",
x"00A9",
x"00A8",
x"00A8",
x"00A9",
x"00A7",
x"00A6",
x"00A8",
x"00A7",
x"00A6",
x"00A8",
x"00A7",
x"00A5",
x"00A5",
x"00A6",
x"00A3",
x"00A7",
x"00A5",
x"00A5",
x"00A5",
x"00A6",
x"00A5",
x"00A6",
x"00A7",
x"00A5",
x"00A5",
x"00A7",
x"00A7",
x"00A5",
x"00A5",
x"00A6",
x"00A5",
x"00A6",
x"00A4",
x"00A4",
x"00A5",
x"00A5",
x"00A3",
x"00A6",
x"00A7",
x"00A6",
x"00A7",
x"00A6",
x"00A5",
x"00A5",
x"00A5",
x"00A5",
x"00A7",
x"00A7",
x"00A6",
x"00A6",
x"00A6",
x"00A6",
x"00A6",
x"00A8",
x"00A7",
x"00A6",
x"00A6",
x"00A6",
x"00B2",
x"00A3",
x"009D",
x"00A1",
x"008C",
x"006A",
x"0070",
x"006A",
x"0049",
x"0029",
x"000F",
x"0057",
x"009B",
x"009E",
x"009D",
x"0090",
x"0085",
x"0088",
x"0084",
x"0084",
x"008F",
x"008A",
x"007D",
x"008F",
x"008D",
x"0087",
x"0082",
x"0087",
x"0092",
x"008A",
x"0077",
x"007E",
x"008A",
x"0095",
x"0081",
x"007E",
x"0081",
x"007F",
x"008B",
x"0080",
x"0089",
x"007D",
x"0072",
x"0083",
x"0085",
x"007E",
x"0082",
x"0083",
x"0083",
x"0084",
x"0078",
x"0097",
x"0000",
x"0000",
x"0000",
x"0000",
x"00AA",
x"00AA",
x"00A9",
x"00A7",
x"00A9",
x"00AA",
x"00A9",
x"00A8",
x"00AA",
x"00AA",
x"00A9",
x"00AD",
x"00AA",
x"00AB",
x"00AC",
x"00A9",
x"00A7",
x"00A8",
x"00AA",
x"00A7",
x"00A8",
x"00A7",
x"00A7",
x"00A7",
x"00A7",
x"00A6",
x"00A5",
x"00A8",
x"00A6",
x"00A4",
x"00A4",
x"00A5",
x"00A4",
x"00A5",
x"00A5",
x"00A3",
x"00A3",
x"00A5",
x"00A4",
x"00A5",
x"00A7",
x"00A4",
x"00A3",
x"00A6",
x"00A6",
x"00A5",
x"00A7",
x"00A6",
x"00A5",
x"00A5",
x"00A6",
x"00A3",
x"00A0",
x"00A4",
x"00A4",
x"00A6",
x"00A5",
x"00A4",
x"00A5",
x"00A5",
x"00A4",
x"00A4",
x"00A5",
x"00A6",
x"00A6",
x"00A7",
x"00A7",
x"00A6",
x"00A6",
x"00A5",
x"00A6",
x"00A8",
x"00A7",
x"00A6",
x"00A6",
x"00A6",
x"00B2",
x"00A3",
x"009A",
x"0089",
x"007E",
x"0043",
x"004A",
x"0047",
x"002E",
x"001A",
x"000D",
x"0059",
x"009B",
x"009C",
x"009D",
x"0092",
x"0082",
x"008A",
x"0080",
x"007E",
x"008C",
x"008B",
x"007B",
x"0092",
x"0090",
x"0083",
x"0081",
x"008B",
x"00A1",
x"0087",
x"007A",
x"0088",
x"0087",
x"0099",
x"008C",
x"0076",
x"007F",
x"0085",
x"008C",
x"0086",
x"008F",
x"0085",
x"006F",
x"0078",
x"0077",
x"008A",
x"006F",
x"0083",
x"007E",
x"0089",
x"008B",
x"009F",
x"0000",
x"0000",
x"0000",
x"0000",
x"00A9",
x"00AA",
x"00A8",
x"00A6",
x"00A7",
x"00A9",
x"00A9",
x"00A8",
x"00A9",
x"00AB",
x"00AB",
x"00AB",
x"00AA",
x"00AA",
x"00AB",
x"00A9",
x"00A8",
x"00A9",
x"00AA",
x"00A9",
x"00A8",
x"00A7",
x"00A7",
x"00A7",
x"00A7",
x"00A5",
x"00A5",
x"00A7",
x"00A7",
x"00A4",
x"00A4",
x"00A4",
x"00A3",
x"00A5",
x"00A5",
x"00A3",
x"00A3",
x"00A4",
x"00A3",
x"00A4",
x"00A6",
x"00A5",
x"00A4",
x"00A5",
x"00A4",
x"00A4",
x"00A5",
x"00A5",
x"00A3",
x"00A3",
x"00A3",
x"00A3",
x"00A5",
x"00A4",
x"00A4",
x"00A6",
x"00A5",
x"00A3",
x"00A4",
x"00A4",
x"00A4",
x"00A4",
x"00A4",
x"00A6",
x"00A6",
x"00A7",
x"00A6",
x"00A4",
x"00A6",
x"00A6",
x"00A5",
x"00A6",
x"00A5",
x"00A4",
x"00A6",
x"00A5",
x"00B3",
x"00A1",
x"0090",
x"007C",
x"0076",
x"0045",
x"0045",
x"004A",
x"0038",
x"001F",
x"0011",
x"005B",
x"009A",
x"009B",
x"009D",
x"008F",
x"0080",
x"0088",
x"0080",
x"007D",
x"008B",
x"0088",
x"0074",
x"008D",
x"0091",
x"0081",
x"007E",
x"0088",
x"009C",
x"0088",
x"0071",
x"0082",
x"0083",
x"0092",
x"0089",
x"0080",
x"0081",
x"0080",
x"0087",
x"007A",
x"0083",
x"0079",
x"0072",
x"0081",
x"008A",
x"009A",
x"0075",
x"0087",
x"0097",
x"0084",
x"0081",
x"0098",
x"0000",
x"0000",
x"0000",
x"0000",
x"00AA",
x"00AA",
x"00A9",
x"00A8",
x"00A8",
x"00A9",
x"00AA",
x"00A9",
x"00AB",
x"00AB",
x"00AA",
x"00AD",
x"00AC",
x"00AA",
x"00A9",
x"00A8",
x"00A9",
x"00AA",
x"00AB",
x"00A8",
x"00A8",
x"00A8",
x"00A7",
x"00A7",
x"00A8",
x"00A5",
x"00A6",
x"00A7",
x"00A7",
x"00A5",
x"00A7",
x"00A4",
x"00A2",
x"00A5",
x"00A4",
x"00A2",
x"00A3",
x"00A3",
x"00A2",
x"00A2",
x"00A4",
x"00A4",
x"00A3",
x"00A4",
x"00A4",
x"00A4",
x"00A3",
x"00A3",
x"00A2",
x"00A2",
x"00A2",
x"00A2",
x"00A4",
x"00A3",
x"00A4",
x"00A4",
x"00A5",
x"00A4",
x"00A5",
x"00A3",
x"00A3",
x"00A3",
x"00A4",
x"00A6",
x"00A7",
x"00A6",
x"00A4",
x"00A3",
x"00A5",
x"00A6",
x"00A4",
x"00A4",
x"00A5",
x"00A4",
x"00A4",
x"00A7",
x"00B5",
x"00A4",
x"0092",
x"0068",
x"005E",
x"005A",
x"0045",
x"004C",
x"0047",
x"0024",
x"0014",
x"0060",
x"0099",
x"009E",
x"009C",
x"008C",
x"007B",
x"0086",
x"007F",
x"007D",
x"0089",
x"0086",
x"0074",
x"0089",
x"0090",
x"007E",
x"0077",
x"008A",
x"009B",
x"008A",
x"006E",
x"0083",
x"0087",
x"008E",
x"008E",
x"008F",
x"0086",
x"0085",
x"0088",
x"007E",
x"008E",
x"0085",
x"007E",
x"0083",
x"0091",
x"0086",
x"0081",
x"0086",
x"007D",
x"007A",
x"007F",
x"0083",
x"0000",
x"0000",
x"0000",
x"0000",
x"00AA",
x"00AA",
x"00A8",
x"00A6",
x"00A7",
x"00A9",
x"00A9",
x"00AA",
x"00AC",
x"00AB",
x"00AB",
x"00AD",
x"00AB",
x"00A9",
x"00AB",
x"00A9",
x"00A8",
x"00AA",
x"00AA",
x"00A7",
x"00A8",
x"00A7",
x"00A6",
x"00A7",
x"00A7",
x"00A6",
x"00A7",
x"00A7",
x"00A7",
x"00A5",
x"00A5",
x"00A4",
x"00A3",
x"00A5",
x"00A3",
x"00A1",
x"00A2",
x"00A4",
x"00A1",
x"00A1",
x"00A4",
x"00A4",
x"00A2",
x"00A5",
x"00A5",
x"00A2",
x"00A2",
x"00A3",
x"00A2",
x"00A1",
x"00A1",
x"00A0",
x"00A2",
x"00A2",
x"00A3",
x"00A4",
x"00A5",
x"00A4",
x"00A5",
x"00A3",
x"00A3",
x"00A4",
x"00A5",
x"00A5",
x"00A5",
x"00A5",
x"00A5",
x"00A4",
x"00A5",
x"00A5",
x"00A4",
x"00A5",
x"00A3",
x"00A4",
x"00A5",
x"00A7",
x"00B3",
x"00A2",
x"009C",
x"0077",
x"0070",
x"006D",
x"0059",
x"004C",
x"0043",
x"002E",
x"0023",
x"0066",
x"0097",
x"009D",
x"009C",
x"008F",
x"007E",
x"0080",
x"007A",
x"007F",
x"008D",
x"008B",
x"007A",
x"0089",
x"0092",
x"0086",
x"0082",
x"008D",
x"0098",
x"0096",
x"0078",
x"0075",
x"0087",
x"0092",
x"008D",
x"008A",
x"0082",
x"0082",
x"0087",
x"007F",
x"0090",
x"0084",
x"0093",
x"0096",
x"0091",
x"0082",
x"007A",
x"008D",
x"0081",
x"007B",
x"0083",
x"0082",
x"0000",
x"0000",
x"0000",
x"0000",
x"00AB",
x"00AB",
x"00A8",
x"00A7",
x"00A7",
x"00A8",
x"00A9",
x"00AA",
x"00AB",
x"00AA",
x"00AB",
x"00AD",
x"00A9",
x"00A7",
x"00A9",
x"00A9",
x"00A8",
x"00AB",
x"00AA",
x"00A8",
x"00A8",
x"00A6",
x"00A5",
x"00A7",
x"00A8",
x"00A4",
x"00A4",
x"00A7",
x"00A7",
x"00A4",
x"00A4",
x"00A4",
x"00A4",
x"00A4",
x"00A3",
x"00A2",
x"00A4",
x"00A3",
x"00A1",
x"00A1",
x"00A4",
x"00A3",
x"00A2",
x"00A3",
x"00A3",
x"00A1",
x"00A2",
x"00A3",
x"00A2",
x"00A1",
x"00A0",
x"00A1",
x"00A1",
x"00A1",
x"00A0",
x"00A2",
x"00A2",
x"00A2",
x"00A3",
x"00A3",
x"00A2",
x"00A3",
x"00A3",
x"00A3",
x"00A6",
x"00A5",
x"00A4",
x"00A4",
x"00A4",
x"00A6",
x"00A4",
x"00A4",
x"00A3",
x"00A3",
x"00A5",
x"00A9",
x"00B5",
x"009E",
x"00A4",
x"0095",
x"0084",
x"0071",
x"006F",
x"005F",
x"003F",
x"0029",
x"001F",
x"0067",
x"0099",
x"009C",
x"009A",
x"008E",
x"007F",
x"0086",
x"007C",
x"007A",
x"008A",
x"0087",
x"007C",
x"008D",
x"008B",
x"0089",
x"008C",
x"0092",
x"0096",
x"008A",
x"0070",
x"0079",
x"0083",
x"0086",
x"008A",
x"0080",
x"0076",
x"0092",
x"008E",
x"007C",
x"0090",
x"0092",
x"008E",
x"0086",
x"0082",
x"008B",
x"007E",
x"0086",
x"0090",
x"0079",
x"0079",
x"0078",
x"0000",
x"0000",
x"0000",
x"0000",
x"00AB",
x"00AB",
x"00A7",
x"00A6",
x"00A6",
x"00A8",
x"00A8",
x"00A6",
x"00A8",
x"00A8",
x"00AB",
x"00AD",
x"00AA",
x"00A8",
x"00A9",
x"00A8",
x"00A7",
x"00A8",
x"00A9",
x"00A7",
x"00A7",
x"00A7",
x"00A6",
x"00A7",
x"00A7",
x"00A7",
x"00A4",
x"00A6",
x"00A5",
x"00A3",
x"00A3",
x"00A2",
x"00A0",
x"00A3",
x"00A3",
x"00A2",
x"00A3",
x"00A3",
x"00A2",
x"00A1",
x"00A3",
x"00A2",
x"00A1",
x"00A2",
x"00A2",
x"00A1",
x"00A2",
x"00A3",
x"00A0",
x"009F",
x"00A0",
x"009F",
x"00A0",
x"009F",
x"009F",
x"00A1",
x"00A0",
x"00A1",
x"00A1",
x"00A1",
x"00A1",
x"00A2",
x"00A1",
x"00A2",
x"00A4",
x"00A2",
x"00A3",
x"00A3",
x"00A4",
x"00A4",
x"00A2",
x"00A3",
x"00A3",
x"00A3",
x"00A4",
x"00A6",
x"00B4",
x"009C",
x"009A",
x"0064",
x"006E",
x"0065",
x"005A",
x"0052",
x"0034",
x"0026",
x"001C",
x"0061",
x"0099",
x"009B",
x"009A",
x"008E",
x"0081",
x"0084",
x"0073",
x"0077",
x"0087",
x"007E",
x"0078",
x"008F",
x"008A",
x"0088",
x"0081",
x"0087",
x"009D",
x"0090",
x"005F",
x"0078",
x"0081",
x"0087",
x"008E",
x"007E",
x"0080",
x"0090",
x"008F",
x"0081",
x"0095",
x"008F",
x"0095",
x"0088",
x"007F",
x"007C",
x"007D",
x"0083",
x"0094",
x"007D",
x"007D",
x"0091",
x"0000",
x"0000",
x"0000",
x"0000",
x"00A9",
x"00A9",
x"00A6",
x"00A5",
x"00A6",
x"00A8",
x"00A8",
x"00A6",
x"00A8",
x"00A9",
x"00A9",
x"00AC",
x"00A9",
x"00A8",
x"00A9",
x"00A8",
x"00A7",
x"00A8",
x"00A8",
x"00A6",
x"00A6",
x"00A6",
x"00A5",
x"00A3",
x"00A6",
x"00A5",
x"00A2",
x"00A4",
x"00A5",
x"00A3",
x"00A4",
x"00A3",
x"00A1",
x"00A1",
x"00A2",
x"00A2",
x"00A2",
x"00A3",
x"00A2",
x"00A3",
x"00A3",
x"00A3",
x"00A1",
x"00A2",
x"00A2",
x"00A2",
x"00A1",
x"00A2",
x"009F",
x"009F",
x"009F",
x"009E",
x"009E",
x"009F",
x"009E",
x"00A0",
x"009E",
x"00A0",
x"00A0",
x"00A0",
x"00A2",
x"00A1",
x"00A2",
x"00A1",
x"00A3",
x"00A2",
x"00A1",
x"00A2",
x"00A3",
x"00A3",
x"00A2",
x"00A2",
x"00A3",
x"00A3",
x"00A3",
x"00A5",
x"00B3",
x"009C",
x"00A7",
x"0082",
x"006A",
x"0065",
x"005D",
x"004F",
x"003A",
x"002A",
x"001F",
x"0060",
x"0098",
x"0099",
x"0098",
x"008E",
x"0080",
x"0082",
x"0078",
x"007B",
x"0087",
x"0081",
x"007E",
x"0091",
x"008D",
x"008B",
x"0087",
x"0082",
x"0096",
x"0096",
x"0056",
x"006C",
x"0086",
x"008B",
x"008B",
x"007D",
x"008A",
x"008A",
x"0099",
x"007D",
x"0082",
x"0088",
x"0092",
x"0085",
x"008A",
x"0082",
x"0081",
x"0095",
x"0094",
x"0070",
x"008C",
x"0095",
x"0000",
x"0000",
x"0000",
x"0000",
x"00A8",
x"00A7",
x"00A8",
x"00A6",
x"00A5",
x"00A8",
x"00A7",
x"00A7",
x"00A8",
x"00A9",
x"00A8",
x"00AB",
x"00A9",
x"00A8",
x"00A9",
x"00A7",
x"00A7",
x"00A7",
x"00A7",
x"00A6",
x"00A6",
x"00A8",
x"00A6",
x"00A6",
x"00A7",
x"00A3",
x"00A2",
x"00A4",
x"00A4",
x"00A2",
x"00A3",
x"00A2",
x"00A0",
x"00A2",
x"00A3",
x"00A1",
x"00A1",
x"00A2",
x"00A2",
x"00A1",
x"00A3",
x"00A2",
x"00A0",
x"00A1",
x"00A1",
x"00A0",
x"00A0",
x"00A2",
x"009F",
x"009F",
x"009F",
x"009E",
x"009D",
x"009E",
x"009E",
x"00A0",
x"00A0",
x"009E",
x"009F",
x"00A0",
x"00A0",
x"00A2",
x"00A3",
x"00A2",
x"00A2",
x"00A2",
x"00A2",
x"00A2",
x"00A2",
x"00A4",
x"00A4",
x"00A4",
x"00A4",
x"00A2",
x"00A3",
x"00A3",
x"00B1",
x"009B",
x"009E",
x"006F",
x"005A",
x"005F",
x"005E",
x"0056",
x"0040",
x"0027",
x"001D",
x"0061",
x"009A",
x"0099",
x"0097",
x"008C",
x"0083",
x"007F",
x"007B",
x"007F",
x"008A",
x"008A",
x"007F",
x"0093",
x"0091",
x"008F",
x"0084",
x"0086",
x"0096",
x"0091",
x"005C",
x"006C",
x"0084",
x"0089",
x"0085",
x"007E",
x"0081",
x"007F",
x"0090",
x"0077",
x"0075",
x"008C",
x"008F",
x"0079",
x"008E",
x"0087",
x"0085",
x"0088",
x"0083",
x"0076",
x"008D",
x"008D",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000");

  signal read_en_int, write_en_int: std_logic;
  signal address_int: std_logic_vector(14 downto 0);
  begin
    main : process(clock)
      begin
        if rising_edge(clock) then
          read_en_int <= rden;
          address_int <= address;
          write_en_int <= wren;
          -- int_data <= data;
          if write_en_int = '1' then
            memory(to_integer(unsigned(address))) <= data;
          end if;
        end if;
      end process;
      q <= memory(to_integer(unsigned(address_int)));-- when read_en_int = '1' else (others => 'Z');
end architecture;
